module tokenizer

const (
	char_ref = {
		'Aacute;':                          [rune(0x000C1)]
		'Aacute':                           [rune(0x000C1)]
		'aacute;':                          [rune(0x000E1)]
		'aacute':                           [rune(0x000E1)]
		'Abreve;':                          [rune(0x00102)]
		'abreve;':                          [rune(0x00103)]
		'ac;':                              [rune(0x0223E)]
		'acd;':                             [rune(0x0223F)]
		'acE;':                             [rune(0x0223E), 0x00333]
		'Acirc;':                           [rune(0x000C2)]
		'Acirc':                            [rune(0x000C2)]
		'acirc;':                           [rune(0x000E2)]
		'acirc':                            [rune(0x000E2)]
		'acute;':                           [rune(0x000B4)]
		'acute':                            [rune(0x000B4)]
		'Acy;':                             [rune(0x00410)]
		'acy;':                             [rune(0x00430)]
		'AElig;':                           [rune(0x000C6)]
		'AElig':                            [rune(0x000C6)]
		'aelig;':                           [rune(0x000E6)]
		'aelig':                            [rune(0x000E6)]
		'af;':                              [rune(0x02061)]
		'Afr;':                             [rune(0x1D504)]
		'afr;':                             [rune(0x1D51E)]
		'Agrave;':                          [rune(0x000C0)]
		'Agrave':                           [rune(0x000C0)]
		'agrave;':                          [rune(0x000E0)]
		'agrave':                           [rune(0x000E0)]
		'alefsym;':                         [rune(0x02135)]
		'aleph;':                           [rune(0x02135)]
		'Alpha;':                           [rune(0x00391)]
		'alpha;':                           [rune(0x003B1)]
		'Amacr;':                           [rune(0x00100)]
		'amacr;':                           [rune(0x00101)]
		'amalg;':                           [rune(0x02A3F)]
		'AMP;':                             [rune(0x00026)]
		'AMP':                              [rune(0x00026)]
		'amp;':                             [rune(0x00026)]
		'amp':                              [rune(0x00026)]
		'And;':                             [rune(0x02A53)]
		'and;':                             [rune(0x02227)]
		'andand;':                          [rune(0x02A55)]
		'andd;':                            [rune(0x02A5C)]
		'andslope;':                        [rune(0x02A58)]
		'andv;':                            [rune(0x02A5A)]
		'ang;':                             [rune(0x02220)]
		'ange;':                            [rune(0x029A4)]
		'angle;':                           [rune(0x02220)]
		'angmsd;':                          [rune(0x02221)]
		'angmsdaa;':                        [rune(0x029A8)]
		'angmsdab;':                        [rune(0x029A9)]
		'angmsdac;':                        [rune(0x029AA)]
		'angmsdad;':                        [rune(0x029AB)]
		'angmsdae;':                        [rune(0x029AC)]
		'angmsdaf;':                        [rune(0x029AD)]
		'angmsdag;':                        [rune(0x029AE)]
		'angmsdah;':                        [rune(0x029AF)]
		'angrt;':                           [rune(0x0221F)]
		'angrtvb;':                         [rune(0x022BE)]
		'angrtvbd;':                        [rune(0x0299D)]
		'angsph;':                          [rune(0x02222)]
		'angst;':                           [rune(0x000C5)]
		'angzarr;':                         [rune(0x0237C)]
		'Aogon;':                           [rune(0x00104)]
		'aogon;':                           [rune(0x00105)]
		'Aopf;':                            [rune(0x1D538)]
		'aopf;':                            [rune(0x1D552)]
		'ap;':                              [rune(0x02248)]
		'apacir;':                          [rune(0x02A6F)]
		'apE;':                             [rune(0x02A70)]
		'ape;':                             [rune(0x0224A)]
		'apid;':                            [rune(0x0224B)]
		'apos;':                            [rune(0x00027)]
		'ApplyFunction;':                   [rune(0x02061)]
		'approx;':                          [rune(0x02248)]
		'approxeq;':                        [rune(0x0224A)]
		'Aring;':                           [rune(0x000C5)]
		'Aring':                            [rune(0x000C5)]
		'aring;':                           [rune(0x000E5)]
		'aring':                            [rune(0x000E5)]
		'Ascr;':                            [rune(0x1D49C)]
		'ascr;':                            [rune(0x1D4B6)]
		'Assign;':                          [rune(0x02254)]
		'ast;':                             [rune(0x0002A)]
		'asymp;':                           [rune(0x02248)]
		'asympeq;':                         [rune(0x0224D)]
		'Atilde;':                          [rune(0x000C3)]
		'Atilde':                           [rune(0x000C3)]
		'atilde;':                          [rune(0x000E3)]
		'atilde':                           [rune(0x000E3)]
		'Auml;':                            [rune(0x000C4)]
		'Auml':                             [rune(0x000C4)]
		'auml;':                            [rune(0x000E4)]
		'auml':                             [rune(0x000E4)]
		'awconint;':                        [rune(0x02233)]
		'awint;':                           [rune(0x02A11)]
		'backcong;':                        [rune(0x0224C)]
		'backepsilon;':                     [rune(0x003F6)]
		'backprime;':                       [rune(0x02035)]
		'backsim;':                         [rune(0x0223D)]
		'backsimeq;':                       [rune(0x022CD)]
		'Backslash;':                       [rune(0x02216)]
		'Barv;':                            [rune(0x02AE7)]
		'barvee;':                          [rune(0x022BD)]
		'Barwed;':                          [rune(0x02306)]
		'barwed;':                          [rune(0x02305)]
		'barwedge;':                        [rune(0x02305)]
		'bbrk;':                            [rune(0x023B5)]
		'bbrktbrk;':                        [rune(0x023B6)]
		'bcong;':                           [rune(0x0224C)]
		'Bcy;':                             [rune(0x00411)]
		'bcy;':                             [rune(0x00431)]
		'bdquo;':                           [rune(0x0201E)]
		'becaus;':                          [rune(0x02235)]
		'Because;':                         [rune(0x02235)]
		'because;':                         [rune(0x02235)]
		'bemptyv;':                         [rune(0x029B0)]
		'bepsi;':                           [rune(0x003F6)]
		'bernou;':                          [rune(0x0212C)]
		'Bernoullis;':                      [rune(0x0212C)]
		'Beta;':                            [rune(0x00392)]
		'beta;':                            [rune(0x003B2)]
		'beth;':                            [rune(0x02136)]
		'between;':                         [rune(0x0226C)]
		'Bfr;':                             [rune(0x1D505)]
		'bfr;':                             [rune(0x1D51F)]
		'bigcap;':                          [rune(0x022C2)]
		'bigcirc;':                         [rune(0x025EF)]
		'bigcup;':                          [rune(0x022C3)]
		'bigodot;':                         [rune(0x02A00)]
		'bigoplus;':                        [rune(0x02A01)]
		'bigotimes;':                       [rune(0x02A02)]
		'bigsqcup;':                        [rune(0x02A06)]
		'bigstar;':                         [rune(0x02605)]
		'bigtriangledown;':                 [rune(0x025BD)]
		'bigtriangleup;':                   [rune(0x025B3)]
		'biguplus;':                        [rune(0x02A04)]
		'bigvee;':                          [rune(0x022C1)]
		'bigwedge;':                        [rune(0x022C0)]
		'bkarow;':                          [rune(0x0290D)]
		'blacklozenge;':                    [rune(0x029EB)]
		'blacksquare;':                     [rune(0x025AA)]
		'blacktriangle;':                   [rune(0x025B4)]
		'blacktriangledown;':               [rune(0x025BE)]
		'blacktriangleleft;':               [rune(0x025C2)]
		'blacktriangleright;':              [rune(0x025B8)]
		'blank;':                           [rune(0x02423)]
		'blk12;':                           [rune(0x02592)]
		'blk14;':                           [rune(0x02591)]
		'blk34;':                           [rune(0x02593)]
		'block;':                           [rune(0x02588)]
		'bne;':                             [rune(0x0003D), 0x020E5]
		'bnequiv;':                         [rune(0x02261), 0x020E5]
		'bNot;':                            [rune(0x02AED)]
		'bnot;':                            [rune(0x02310)]
		'Bopf;':                            [rune(0x1D539)]
		'bopf;':                            [rune(0x1D553)]
		'bot;':                             [rune(0x022A5)]
		'bottom;':                          [rune(0x022A5)]
		'bowtie;':                          [rune(0x022C8)]
		'boxbox;':                          [rune(0x029C9)]
		'boxDL;':                           [rune(0x02557)]
		'boxDl;':                           [rune(0x02556)]
		'boxdL;':                           [rune(0x02555)]
		'boxdl;':                           [rune(0x02510)]
		'boxDR;':                           [rune(0x02554)]
		'boxDr;':                           [rune(0x02553)]
		'boxdR;':                           [rune(0x02552)]
		'boxdr;':                           [rune(0x0250C)]
		'boxH;':                            [rune(0x02550)]
		'boxh;':                            [rune(0x02500)]
		'boxHD;':                           [rune(0x02566)]
		'boxHd;':                           [rune(0x02564)]
		'boxhD;':                           [rune(0x02565)]
		'boxhd;':                           [rune(0x0252C)]
		'boxHU;':                           [rune(0x02569)]
		'boxHu;':                           [rune(0x02567)]
		'boxhU;':                           [rune(0x02568)]
		'boxhu;':                           [rune(0x02534)]
		'boxminus;':                        [rune(0x0229F)]
		'boxplus;':                         [rune(0x0229E)]
		'boxtimes;':                        [rune(0x022A0)]
		'boxUL;':                           [rune(0x0255D)]
		'boxUl;':                           [rune(0x0255C)]
		'boxuL;':                           [rune(0x0255B)]
		'boxul;':                           [rune(0x02518)]
		'boxUR;':                           [rune(0x0255A)]
		'boxUr;':                           [rune(0x02559)]
		'boxuR;':                           [rune(0x02558)]
		'boxur;':                           [rune(0x02514)]
		'boxV;':                            [rune(0x02551)]
		'boxv;':                            [rune(0x02502)]
		'boxVH;':                           [rune(0x0256C)]
		'boxVh;':                           [rune(0x0256B)]
		'boxvH;':                           [rune(0x0256A)]
		'boxvh;':                           [rune(0x0253C)]
		'boxVL;':                           [rune(0x02563)]
		'boxVl;':                           [rune(0x02562)]
		'boxvL;':                           [rune(0x02561)]
		'boxvl;':                           [rune(0x02524)]
		'boxVR;':                           [rune(0x02560)]
		'boxVr;':                           [rune(0x0255F)]
		'boxvR;':                           [rune(0x0255E)]
		'boxvr;':                           [rune(0x0251C)]
		'bprime;':                          [rune(0x02035)]
		'Breve;':                           [rune(0x002D8)]
		'breve;':                           [rune(0x002D8)]
		'brvbar;':                          [rune(0x000A6)]
		'brvbar':                           [rune(0x000A6)]
		'Bscr;':                            [rune(0x0212C)]
		'bscr;':                            [rune(0x1D4B7)]
		'bsemi;':                           [rune(0x0204F)]
		'bsim;':                            [rune(0x0223D)]
		'bsime;':                           [rune(0x022CD)]
		'bsol;':                            [rune(0x0005C)]
		'bsolb;':                           [rune(0x029C5)]
		'bsolhsub;':                        [rune(0x027C8)]
		'bull;':                            [rune(0x02022)]
		'bullet;':                          [rune(0x02022)]
		'bump;':                            [rune(0x0224E)]
		'bumpE;':                           [rune(0x02AAE)]
		'bumpe;':                           [rune(0x0224F)]
		'Bumpeq;':                          [rune(0x0224E)]
		'bumpeq;':                          [rune(0x0224F)]
		'Cacute;':                          [rune(0x00106)]
		'cacute;':                          [rune(0x00107)]
		'Cap;':                             [rune(0x022D2)]
		'cap;':                             [rune(0x02229)]
		'capand;':                          [rune(0x02A44)]
		'capbrcup;':                        [rune(0x02A49)]
		'capcap;':                          [rune(0x02A4B)]
		'capcup;':                          [rune(0x02A47)]
		'capdot;':                          [rune(0x02A40)]
		'CapitalDifferentialD;':            [rune(0x02145)]
		'caps;':                            [rune(0x02229), 0x0FE00]
		'caret;':                           [rune(0x02041)]
		'caron;':                           [rune(0x002C7)]
		'Cayleys;':                         [rune(0x0212D)]
		'ccaps;':                           [rune(0x02A4D)]
		'Ccaron;':                          [rune(0x0010C)]
		'ccaron;':                          [rune(0x0010D)]
		'Ccedil;':                          [rune(0x000C7)]
		'Ccedil':                           [rune(0x000C7)]
		'ccedil;':                          [rune(0x000E7)]
		'ccedil':                           [rune(0x000E7)]
		'Ccirc;':                           [rune(0x00108)]
		'ccirc;':                           [rune(0x00109)]
		'Cconint;':                         [rune(0x02230)]
		'ccups;':                           [rune(0x02A4C)]
		'ccupssm;':                         [rune(0x02A50)]
		'Cdot;':                            [rune(0x0010A)]
		'cdot;':                            [rune(0x0010B)]
		'cedil;':                           [rune(0x000B8)]
		'cedil':                            [rune(0x000B8)]
		'Cedilla;':                         [rune(0x000B8)]
		'cemptyv;':                         [rune(0x029B2)]
		'cent;':                            [rune(0x000A2)]
		'cent':                             [rune(0x000A2)]
		'CenterDot;':                       [rune(0x000B7)]
		'centerdot;':                       [rune(0x000B7)]
		'Cfr;':                             [rune(0x0212D)]
		'cfr;':                             [rune(0x1D520)]
		'CHcy;':                            [rune(0x00427)]
		'chcy;':                            [rune(0x00447)]
		'check;':                           [rune(0x02713)]
		'checkmark;':                       [rune(0x02713)]
		'Chi;':                             [rune(0x003A7)]
		'chi;':                             [rune(0x003C7)]
		'cir;':                             [rune(0x025CB)]
		'circ;':                            [rune(0x002C6)]
		'circeq;':                          [rune(0x02257)]
		'circlearrowleft;':                 [rune(0x021BA)]
		'circlearrowright;':                [rune(0x021BB)]
		'circledast;':                      [rune(0x0229B)]
		'circledcirc;':                     [rune(0x0229A)]
		'circleddash;':                     [rune(0x0229D)]
		'CircleDot;':                       [rune(0x02299)]
		'circledR;':                        [rune(0x000AE)]
		'circledS;':                        [rune(0x024C8)]
		'CircleMinus;':                     [rune(0x02296)]
		'CirclePlus;':                      [rune(0x02295)]
		'CircleTimes;':                     [rune(0x02297)]
		'cirE;':                            [rune(0x029C3)]
		'cire;':                            [rune(0x02257)]
		'cirfnint;':                        [rune(0x02A10)]
		'cirmid;':                          [rune(0x02AEF)]
		'cirscir;':                         [rune(0x029C2)]
		'ClockwiseContourIntegral;':        [rune(0x02232)]
		'CloseCurlyDoubleQuote;':           [rune(0x0201D)]
		'CloseCurlyQuote;':                 [rune(0x02019)]
		'clubs;':                           [rune(0x02663)]
		'clubsuit;':                        [rune(0x02663)]
		'Colon;':                           [rune(0x02237)]
		'colon;':                           [rune(0x0003A)]
		'Colone;':                          [rune(0x02A74)]
		'colone;':                          [rune(0x02254)]
		'coloneq;':                         [rune(0x02254)]
		'comma;':                           [rune(0x0002C)]
		'commat;':                          [rune(0x00040)]
		'comp;':                            [rune(0x02201)]
		'compfn;':                          [rune(0x02218)]
		'complement;':                      [rune(0x02201)]
		'complexes;':                       [rune(0x02102)]
		'cong;':                            [rune(0x02245)]
		'congdot;':                         [rune(0x02A6D)]
		'Congruent;':                       [rune(0x02261)]
		'Conint;':                          [rune(0x0222F)]
		'conint;':                          [rune(0x0222E)]
		'ContourIntegral;':                 [rune(0x0222E)]
		'Copf;':                            [rune(0x02102)]
		'copf;':                            [rune(0x1D554)]
		'coprod;':                          [rune(0x02210)]
		'Coproduct;':                       [rune(0x02210)]
		'COPY;':                            [rune(0x000A9)]
		'COPY':                             [rune(0x000A9)]
		'copy;':                            [rune(0x000A9)]
		'copy':                             [rune(0x000A9)]
		'copysr;':                          [rune(0x02117)]
		'CounterClockwiseContourIntegral;': [rune(0x02233)]
		'crarr;':                           [rune(0x021B5)]
		'Cross;':                           [rune(0x02A2F)]
		'cross;':                           [rune(0x02717)]
		'Cscr;':                            [rune(0x1D49E)]
		'cscr;':                            [rune(0x1D4B8)]
		'csub;':                            [rune(0x02ACF)]
		'csube;':                           [rune(0x02AD1)]
		'csup;':                            [rune(0x02AD0)]
		'csupe;':                           [rune(0x02AD2)]
		'ctdot;':                           [rune(0x022EF)]
		'cudarrl;':                         [rune(0x02938)]
		'cudarrr;':                         [rune(0x02935)]
		'cuepr;':                           [rune(0x022DE)]
		'cuesc;':                           [rune(0x022DF)]
		'cularr;':                          [rune(0x021B6)]
		'cularrp;':                         [rune(0x0293D)]
		'Cup;':                             [rune(0x022D3)]
		'cup;':                             [rune(0x0222A)]
		'cupbrcap;':                        [rune(0x02A48)]
		'CupCap;':                          [rune(0x0224D)]
		'cupcap;':                          [rune(0x02A46)]
		'cupcup;':                          [rune(0x02A4A)]
		'cupdot;':                          [rune(0x0228D)]
		'cupor;':                           [rune(0x02A45)]
		'cups;':                            [rune(0x0222A), 0x0FE00]
		'curarr;':                          [rune(0x021B7)]
		'curarrm;':                         [rune(0x0293C)]
		'curlyeqprec;':                     [rune(0x022DE)]
		'curlyeqsucc;':                     [rune(0x022DF)]
		'curlyvee;':                        [rune(0x022CE)]
		'curlywedge;':                      [rune(0x022CF)]
		'curren;':                          [rune(0x000A4)]
		'curren':                           [rune(0x000A4)]
		'curvearrowleft;':                  [rune(0x021B6)]
		'curvearrowright;':                 [rune(0x021B7)]
		'cuvee;':                           [rune(0x022CE)]
		'cuwed;':                           [rune(0x022CF)]
		'cwconint;':                        [rune(0x02232)]
		'cwint;':                           [rune(0x02231)]
		'cylcty;':                          [rune(0x0232D)]
		'Dagger;':                          [rune(0x02021)]
		'dagger;':                          [rune(0x02020)]
		'daleth;':                          [rune(0x02138)]
		'Darr;':                            [rune(0x021A1)]
		'dArr;':                            [rune(0x021D3)]
		'darr;':                            [rune(0x02193)]
		'dash;':                            [rune(0x02010)]
		'Dashv;':                           [rune(0x02AE4)]
		'dashv;':                           [rune(0x022A3)]
		'dbkarow;':                         [rune(0x0290F)]
		'dblac;':                           [rune(0x002DD)]
		'Dcaron;':                          [rune(0x0010E)]
		'dcaron;':                          [rune(0x0010F)]
		'Dcy;':                             [rune(0x00414)]
		'dcy;':                             [rune(0x00434)]
		'DD;':                              [rune(0x02145)]
		'dd;':                              [rune(0x02146)]
		'ddagger;':                         [rune(0x02021)]
		'ddarr;':                           [rune(0x021CA)]
		'DDotrahd;':                        [rune(0x02911)]
		'ddotseq;':                         [rune(0x02A77)]
		'deg;':                             [rune(0x000B0)]
		'deg':                              [rune(0x000B0)]
		'Del;':                             [rune(0x02207)]
		'Delta;':                           [rune(0x00394)]
		'delta;':                           [rune(0x003B4)]
		'demptyv;':                         [rune(0x029B1)]
		'dfisht;':                          [rune(0x0297F)]
		'Dfr;':                             [rune(0x1D507)]
		'dfr;':                             [rune(0x1D521)]
		'dHar;':                            [rune(0x02965)]
		'dharl;':                           [rune(0x021C3)]
		'dharr;':                           [rune(0x021C2)]
		'DiacriticalAcute;':                [rune(0x000B4)]
		'DiacriticalDot;':                  [rune(0x002D9)]
		'DiacriticalDoubleAcute;':          [rune(0x002DD)]
		'DiacriticalGrave;':                [rune(0x00060)]
		'DiacriticalTilde;':                [rune(0x002DC)]
		'diam;':                            [rune(0x022C4)]
		'Diamond;':                         [rune(0x022C4)]
		'diamond;':                         [rune(0x022C4)]
		'diamondsuit;':                     [rune(0x02666)]
		'diams;':                           [rune(0x02666)]
		'die;':                             [rune(0x000A8)]
		'DifferentialD;':                   [rune(0x02146)]
		'digamma;':                         [rune(0x003DD)]
		'disin;':                           [rune(0x022F2)]
		'div;':                             [rune(0x000F7)]
		'divide;':                          [rune(0x000F7)]
		'divide':                           [rune(0x000F7)]
		'divideontimes;':                   [rune(0x022C7)]
		'divonx;':                          [rune(0x022C7)]
		'DJcy;':                            [rune(0x00402)]
		'djcy;':                            [rune(0x00452)]
		'dlcorn;':                          [rune(0x0231E)]
		'dlcrop;':                          [rune(0x0230D)]
		'dollar;':                          [rune(0x00024)]
		'Dopf;':                            [rune(0x1D53B)]
		'dopf;':                            [rune(0x1D555)]
		'Dot;':                             [rune(0x000A8)]
		'dot;':                             [rune(0x002D9)]
		'DotDot;':                          [rune(0x020DC)]
		'doteq;':                           [rune(0x02250)]
		'doteqdot;':                        [rune(0x02251)]
		'DotEqual;':                        [rune(0x02250)]
		'dotminus;':                        [rune(0x02238)]
		'dotplus;':                         [rune(0x02214)]
		'dotsquare;':                       [rune(0x022A1)]
		'doublebarwedge;':                  [rune(0x02306)]
		'DoubleContourIntegral;':           [rune(0x0222F)]
		'DoubleDot;':                       [rune(0x000A8)]
		'DoubleDownArrow;':                 [rune(0x021D3)]
		'DoubleLeftArrow;':                 [rune(0x021D0)]
		'DoubleLeftRightArrow;':            [rune(0x021D4)]
		'DoubleLeftTee;':                   [rune(0x02AE4)]
		'DoubleLongLeftArrow;':             [rune(0x027F8)]
		'DoubleLongLeftRightArrow;':        [rune(0x027FA)]
		'DoubleLongRightArrow;':            [rune(0x027F9)]
		'DoubleRightArrow;':                [rune(0x021D2)]
		'DoubleRightTee;':                  [rune(0x022A8)]
		'DoubleUpArrow;':                   [rune(0x021D1)]
		'DoubleUpDownArrow;':               [rune(0x021D5)]
		'DoubleVerticalBar;':               [rune(0x02225)]
		'DownArrow;':                       [rune(0x02193)]
		'Downarrow;':                       [rune(0x021D3)]
		'downarrow;':                       [rune(0x02193)]
		'DownArrowBar;':                    [rune(0x02913)]
		'DownArrowUpArrow;':                [rune(0x021F5)]
		'DownBreve;':                       [rune(0x00311)]
		'downdownarrows;':                  [rune(0x021CA)]
		'downharpoonleft;':                 [rune(0x021C3)]
		'downharpoonright;':                [rune(0x021C2)]
		'DownLeftRightVector;':             [rune(0x02950)]
		'DownLeftTeeVector;':               [rune(0x0295E)]
		'DownLeftVector;':                  [rune(0x021BD)]
		'DownLeftVectorBar;':               [rune(0x02956)]
		'DownRightTeeVector;':              [rune(0x0295F)]
		'DownRightVector;':                 [rune(0x021C1)]
		'DownRightVectorBar;':              [rune(0x02957)]
		'DownTee;':                         [rune(0x022A4)]
		'DownTeeArrow;':                    [rune(0x021A7)]
		'drbkarow;':                        [rune(0x02910)]
		'drcorn;':                          [rune(0x0231F)]
		'drcrop;':                          [rune(0x0230C)]
		'Dscr;':                            [rune(0x1D49F)]
		'dscr;':                            [rune(0x1D4B9)]
		'DScy;':                            [rune(0x00405)]
		'dscy;':                            [rune(0x00455)]
		'dsol;':                            [rune(0x029F6)]
		'Dstrok;':                          [rune(0x00110)]
		'dstrok;':                          [rune(0x00111)]
		'dtdot;':                           [rune(0x022F1)]
		'dtri;':                            [rune(0x025BF)]
		'dtrif;':                           [rune(0x025BE)]
		'duarr;':                           [rune(0x021F5)]
		'duhar;':                           [rune(0x0296F)]
		'dwangle;':                         [rune(0x029A6)]
		'DZcy;':                            [rune(0x0040F)]
		'dzcy;':                            [rune(0x0045F)]
		'dzigrarr;':                        [rune(0x027FF)]
		'Eacute;':                          [rune(0x000C9)]
		'Eacute':                           [rune(0x000C9)]
		'eacute;':                          [rune(0x000E9)]
		'eacute':                           [rune(0x000E9)]
		'easter;':                          [rune(0x02A6E)]
		'Ecaron;':                          [rune(0x0011A)]
		'ecaron;':                          [rune(0x0011B)]
		'ecir;':                            [rune(0x02256)]
		'Ecirc;':                           [rune(0x000CA)]
		'Ecirc':                            [rune(0x000CA)]
		'ecirc;':                           [rune(0x000EA)]
		'ecirc':                            [rune(0x000EA)]
		'ecolon;':                          [rune(0x02255)]
		'Ecy;':                             [rune(0x0042D)]
		'ecy;':                             [rune(0x0044D)]
		'eDDot;':                           [rune(0x02A77)]
		'Edot;':                            [rune(0x00116)]
		'eDot;':                            [rune(0x02251)]
		'edot;':                            [rune(0x00117)]
		'ee;':                              [rune(0x02147)]
		'efDot;':                           [rune(0x02252)]
		'Efr;':                             [rune(0x1D508)]
		'efr;':                             [rune(0x1D522)]
		'eg;':                              [rune(0x02A9A)]
		'Egrave;':                          [rune(0x000C8)]
		'Egrave':                           [rune(0x000C8)]
		'egrave;':                          [rune(0x000E8)]
		'egrave':                           [rune(0x000E8)]
		'egs;':                             [rune(0x02A96)]
		'egsdot;':                          [rune(0x02A98)]
		'el;':                              [rune(0x02A99)]
		'Element;':                         [rune(0x02208)]
		'elinters;':                        [rune(0x023E7)]
		'ell;':                             [rune(0x02113)]
		'els;':                             [rune(0x02A95)]
		'elsdot;':                          [rune(0x02A97)]
		'Emacr;':                           [rune(0x00112)]
		'emacr;':                           [rune(0x00113)]
		'empty;':                           [rune(0x02205)]
		'emptyset;':                        [rune(0x02205)]
		'EmptySmallSquare;':                [rune(0x025FB)]
		'emptyv;':                          [rune(0x02205)]
		'EmptyVerySmallSquare;':            [rune(0x025AB)]
		'emsp;':                            [rune(0x02003)]
		'emsp13;':                          [rune(0x02004)]
		'emsp14;':                          [rune(0x02005)]
		'ENG;':                             [rune(0x0014A)]
		'eng;':                             [rune(0x0014B)]
		'ensp;':                            [rune(0x02002)]
		'Eogon;':                           [rune(0x00118)]
		'eogon;':                           [rune(0x00119)]
		'Eopf;':                            [rune(0x1D53C)]
		'eopf;':                            [rune(0x1D556)]
		'epar;':                            [rune(0x022D5)]
		'eparsl;':                          [rune(0x029E3)]
		'eplus;':                           [rune(0x02A71)]
		'epsi;':                            [rune(0x003B5)]
		'Epsilon;':                         [rune(0x00395)]
		'epsilon;':                         [rune(0x003B5)]
		'epsiv;':                           [rune(0x003F5)]
		'eqcirc;':                          [rune(0x02256)]
		'eqcolon;':                         [rune(0x02255)]
		'eqsim;':                           [rune(0x02242)]
		'eqslantgtr;':                      [rune(0x02A96)]
		'eqslantless;':                     [rune(0x02A95)]
		'Equal;':                           [rune(0x02A75)]
		'equals;':                          [rune(0x0003D)]
		'EqualTilde;':                      [rune(0x02242)]
		'equest;':                          [rune(0x0225F)]
		'Equilibrium;':                     [rune(0x021CC)]
		'equiv;':                           [rune(0x02261)]
		'equivDD;':                         [rune(0x02A78)]
		'eqvparsl;':                        [rune(0x029E5)]
		'erarr;':                           [rune(0x02971)]
		'erDot;':                           [rune(0x02253)]
		'Escr;':                            [rune(0x02130)]
		'escr;':                            [rune(0x0212F)]
		'esdot;':                           [rune(0x02250)]
		'Esim;':                            [rune(0x02A73)]
		'esim;':                            [rune(0x02242)]
		'Eta;':                             [rune(0x00397)]
		'eta;':                             [rune(0x003B7)]
		'ETH;':                             [rune(0x000D0)]
		'ETH':                              [rune(0x000D0)]
		'eth;':                             [rune(0x000F0)]
		'eth':                              [rune(0x000F0)]
		'Euml;':                            [rune(0x000CB)]
		'Euml':                             [rune(0x000CB)]
		'euml;':                            [rune(0x000EB)]
		'euml':                             [rune(0x000EB)]
		'euro;':                            [rune(0x020AC)]
		'excl;':                            [rune(0x00021)]
		'exist;':                           [rune(0x02203)]
		'Exists;':                          [rune(0x02203)]
		'expectation;':                     [rune(0x02130)]
		'ExponentialE;':                    [rune(0x02147)]
		'exponentiale;':                    [rune(0x02147)]
		'fallingdotseq;':                   [rune(0x02252)]
		'Fcy;':                             [rune(0x00424)]
		'fcy;':                             [rune(0x00444)]
		'female;':                          [rune(0x02640)]
		'ffilig;':                          [rune(0x0FB03)]
		'fflig;':                           [rune(0x0FB00)]
		'ffllig;':                          [rune(0x0FB04)]
		'Ffr;':                             [rune(0x1D509)]
		'ffr;':                             [rune(0x1D523)]
		'filig;':                           [rune(0x0FB01)]
		'FilledSmallSquare;':               [rune(0x025FC)]
		'FilledVerySmallSquare;':           [rune(0x025AA)]
		'fjlig;':                           [rune(0x00066), 0x0006A]
		'flat;':                            [rune(0x0266D)]
		'fllig;':                           [rune(0x0FB02)]
		'fltns;':                           [rune(0x025B1)]
		'fnof;':                            [rune(0x00192)]
		'Fopf;':                            [rune(0x1D53D)]
		'fopf;':                            [rune(0x1D557)]
		'ForAll;':                          [rune(0x02200)]
		'forall;':                          [rune(0x02200)]
		'fork;':                            [rune(0x022D4)]
		'forkv;':                           [rune(0x02AD9)]
		'Fouriertrf;':                      [rune(0x02131)]
		'fpartint;':                        [rune(0x02A0D)]
		'frac12;':                          [rune(0x000BD)]
		'frac12':                           [rune(0x000BD)]
		'frac13;':                          [rune(0x02153)]
		'frac14;':                          [rune(0x000BC)]
		'frac14':                           [rune(0x000BC)]
		'frac15;':                          [rune(0x02155)]
		'frac16;':                          [rune(0x02159)]
		'frac18;':                          [rune(0x0215B)]
		'frac23;':                          [rune(0x02154)]
		'frac25;':                          [rune(0x02156)]
		'frac34;':                          [rune(0x000BE)]
		'frac34':                           [rune(0x000BE)]
		'frac35;':                          [rune(0x02157)]
		'frac38;':                          [rune(0x0215C)]
		'frac45;':                          [rune(0x02158)]
		'frac56;':                          [rune(0x0215A)]
		'frac58;':                          [rune(0x0215D)]
		'frac78;':                          [rune(0x0215E)]
		'frasl;':                           [rune(0x02044)]
		'frown;':                           [rune(0x02322)]
		'Fscr;':                            [rune(0x02131)]
		'fscr;':                            [rune(0x1D4BB)]
		'gacute;':                          [rune(0x001F5)]
		'Gamma;':                           [rune(0x00393)]
		'gamma;':                           [rune(0x003B3)]
		'Gammad;':                          [rune(0x003DC)]
		'gammad;':                          [rune(0x003DD)]
		'gap;':                             [rune(0x02A86)]
		'Gbreve;':                          [rune(0x0011E)]
		'gbreve;':                          [rune(0x0011F)]
		'Gcedil;':                          [rune(0x00122)]
		'Gcirc;':                           [rune(0x0011C)]
		'gcirc;':                           [rune(0x0011D)]
		'Gcy;':                             [rune(0x00413)]
		'gcy;':                             [rune(0x00433)]
		'Gdot;':                            [rune(0x00120)]
		'gdot;':                            [rune(0x00121)]
		'gE;':                              [rune(0x02267)]
		'ge;':                              [rune(0x02265)]
		'gEl;':                             [rune(0x02A8C)]
		'gel;':                             [rune(0x022DB)]
		'geq;':                             [rune(0x02265)]
		'geqq;':                            [rune(0x02267)]
		'geqslant;':                        [rune(0x02A7E)]
		'ges;':                             [rune(0x02A7E)]
		'gescc;':                           [rune(0x02AA9)]
		'gesdot;':                          [rune(0x02A80)]
		'gesdoto;':                         [rune(0x02A82)]
		'gesdotol;':                        [rune(0x02A84)]
		'gesl;':                            [rune(0x022DB), 0x0FE00]
		'gesles;':                          [rune(0x02A94)]
		'Gfr;':                             [rune(0x1D50A)]
		'gfr;':                             [rune(0x1D524)]
		'Gg;':                              [rune(0x022D9)]
		'gg;':                              [rune(0x0226B)]
		'ggg;':                             [rune(0x022D9)]
		'gimel;':                           [rune(0x02137)]
		'GJcy;':                            [rune(0x00403)]
		'gjcy;':                            [rune(0x00453)]
		'gl;':                              [rune(0x02277)]
		'gla;':                             [rune(0x02AA5)]
		'glE;':                             [rune(0x02A92)]
		'glj;':                             [rune(0x02AA4)]
		'gnap;':                            [rune(0x02A8A)]
		'gnapprox;':                        [rune(0x02A8A)]
		'gnE;':                             [rune(0x02269)]
		'gne;':                             [rune(0x02A88)]
		'gneq;':                            [rune(0x02A88)]
		'gneqq;':                           [rune(0x02269)]
		'gnsim;':                           [rune(0x022E7)]
		'Gopf;':                            [rune(0x1D53E)]
		'gopf;':                            [rune(0x1D558)]
		'grave;':                           [rune(0x00060)]
		'GreaterEqual;':                    [rune(0x02265)]
		'GreaterEqualLess;':                [rune(0x022DB)]
		'GreaterFullEqual;':                [rune(0x02267)]
		'GreaterGreater;':                  [rune(0x02AA2)]
		'GreaterLess;':                     [rune(0x02277)]
		'GreaterSlantEqual;':               [rune(0x02A7E)]
		'GreaterTilde;':                    [rune(0x02273)]
		'Gscr;':                            [rune(0x1D4A2)]
		'gscr;':                            [rune(0x0210A)]
		'gsim;':                            [rune(0x02273)]
		'gsime;':                           [rune(0x02A8E)]
		'gsiml;':                           [rune(0x02A90)]
		'GT;':                              [rune(0x0003E)]
		'GT':                               [rune(0x0003E)]
		'Gt;':                              [rune(0x0226B)]
		'gt;':                              [rune(0x0003E)]
		'gt':                               [rune(0x0003E)]
		'gtcc;':                            [rune(0x02AA7)]
		'gtcir;':                           [rune(0x02A7A)]
		'gtdot;':                           [rune(0x022D7)]
		'gtlPar;':                          [rune(0x02995)]
		'gtquest;':                         [rune(0x02A7C)]
		'gtrapprox;':                       [rune(0x02A86)]
		'gtrarr;':                          [rune(0x02978)]
		'gtrdot;':                          [rune(0x022D7)]
		'gtreqless;':                       [rune(0x022DB)]
		'gtreqqless;':                      [rune(0x02A8C)]
		'gtrless;':                         [rune(0x02277)]
		'gtrsim;':                          [rune(0x02273)]
		'gvertneqq;':                       [rune(0x02269), 0x0FE00]
		'gvnE;':                            [rune(0x02269), 0x0FE00]
		'Hacek;':                           [rune(0x002C7)]
		'hairsp;':                          [rune(0x0200A)]
		'half;':                            [rune(0x000BD)]
		'hamilt;':                          [rune(0x0210B)]
		'HARDcy;':                          [rune(0x0042A)]
		'hardcy;':                          [rune(0x0044A)]
		'hArr;':                            [rune(0x021D4)]
		'harr;':                            [rune(0x02194)]
		'harrcir;':                         [rune(0x02948)]
		'harrw;':                           [rune(0x021AD)]
		'Hat;':                             [rune(0x0005E)]
		'hbar;':                            [rune(0x0210F)]
		'Hcirc;':                           [rune(0x00124)]
		'hcirc;':                           [rune(0x00125)]
		'hearts;':                          [rune(0x02665)]
		'heartsuit;':                       [rune(0x02665)]
		'hellip;':                          [rune(0x02026)]
		'hercon;':                          [rune(0x022B9)]
		'Hfr;':                             [rune(0x0210C)]
		'hfr;':                             [rune(0x1D525)]
		'HilbertSpace;':                    [rune(0x0210B)]
		'hksearow;':                        [rune(0x02925)]
		'hkswarow;':                        [rune(0x02926)]
		'hoarr;':                           [rune(0x021FF)]
		'homtht;':                          [rune(0x0223B)]
		'hookleftarrow;':                   [rune(0x021A9)]
		'hookrightarrow;':                  [rune(0x021AA)]
		'Hopf;':                            [rune(0x0210D)]
		'hopf;':                            [rune(0x1D559)]
		'horbar;':                          [rune(0x02015)]
		'HorizontalLine;':                  [rune(0x02500)]
		'Hscr;':                            [rune(0x0210B)]
		'hscr;':                            [rune(0x1D4BD)]
		'hslash;':                          [rune(0x0210F)]
		'Hstrok;':                          [rune(0x00126)]
		'hstrok;':                          [rune(0x00127)]
		'HumpDownHump;':                    [rune(0x0224E)]
		'HumpEqual;':                       [rune(0x0224F)]
		'hybull;':                          [rune(0x02043)]
		'hyphen;':                          [rune(0x02010)]
		'Iacute;':                          [rune(0x000CD)]
		'Iacute':                           [rune(0x000CD)]
		'iacute;':                          [rune(0x000ED)]
		'iacute':                           [rune(0x000ED)]
		'ic;':                              [rune(0x02063)]
		'Icirc;':                           [rune(0x000CE)]
		'Icirc':                            [rune(0x000CE)]
		'icirc;':                           [rune(0x000EE)]
		'icirc':                            [rune(0x000EE)]
		'Icy;':                             [rune(0x00418)]
		'icy;':                             [rune(0x00438)]
		'Idot;':                            [rune(0x00130)]
		'IEcy;':                            [rune(0x00415)]
		'iecy;':                            [rune(0x00435)]
		'iexcl;':                           [rune(0x000A1)]
		'iexcl':                            [rune(0x000A1)]
		'iff;':                             [rune(0x021D4)]
		'Ifr;':                             [rune(0x02111)]
		'ifr;':                             [rune(0x1D526)]
		'Igrave;':                          [rune(0x000CC)]
		'Igrave':                           [rune(0x000CC)]
		'igrave;':                          [rune(0x000EC)]
		'igrave':                           [rune(0x000EC)]
		'ii;':                              [rune(0x02148)]
		'iiiint;':                          [rune(0x02A0C)]
		'iiint;':                           [rune(0x0222D)]
		'iinfin;':                          [rune(0x029DC)]
		'iiota;':                           [rune(0x02129)]
		'IJlig;':                           [rune(0x00132)]
		'ijlig;':                           [rune(0x00133)]
		'Im;':                              [rune(0x02111)]
		'Imacr;':                           [rune(0x0012A)]
		'imacr;':                           [rune(0x0012B)]
		'image;':                           [rune(0x02111)]
		'ImaginaryI;':                      [rune(0x02148)]
		'imagline;':                        [rune(0x02110)]
		'imagpart;':                        [rune(0x02111)]
		'imath;':                           [rune(0x00131)]
		'imof;':                            [rune(0x022B7)]
		'imped;':                           [rune(0x001B5)]
		'Implies;':                         [rune(0x021D2)]
		'in;':                              [rune(0x02208)]
		'incare;':                          [rune(0x02105)]
		'infin;':                           [rune(0x0221E)]
		'infintie;':                        [rune(0x029DD)]
		'inodot;':                          [rune(0x00131)]
		'Int;':                             [rune(0x0222C)]
		'int;':                             [rune(0x0222B)]
		'intcal;':                          [rune(0x022BA)]
		'integers;':                        [rune(0x02124)]
		'Integral;':                        [rune(0x0222B)]
		'intercal;':                        [rune(0x022BA)]
		'Intersection;':                    [rune(0x022C2)]
		'intlarhk;':                        [rune(0x02A17)]
		'intprod;':                         [rune(0x02A3C)]
		'InvisibleComma;':                  [rune(0x02063)]
		'InvisibleTimes;':                  [rune(0x02062)]
		'IOcy;':                            [rune(0x00401)]
		'iocy;':                            [rune(0x00451)]
		'Iogon;':                           [rune(0x0012E)]
		'iogon;':                           [rune(0x0012F)]
		'Iopf;':                            [rune(0x1D540)]
		'iopf;':                            [rune(0x1D55A)]
		'Iota;':                            [rune(0x00399)]
		'iota;':                            [rune(0x003B9)]
		'iprod;':                           [rune(0x02A3C)]
		'iquest;':                          [rune(0x000BF)]
		'iquest':                           [rune(0x000BF)]
		'Iscr;':                            [rune(0x02110)]
		'iscr;':                            [rune(0x1D4BE)]
		'isin;':                            [rune(0x02208)]
		'isindot;':                         [rune(0x022F5)]
		'isinE;':                           [rune(0x022F9)]
		'isins;':                           [rune(0x022F4)]
		'isinsv;':                          [rune(0x022F3)]
		'isinv;':                           [rune(0x02208)]
		'it;':                              [rune(0x02062)]
		'Itilde;':                          [rune(0x00128)]
		'itilde;':                          [rune(0x00129)]
		'Iukcy;':                           [rune(0x00406)]
		'iukcy;':                           [rune(0x00456)]
		'Iuml;':                            [rune(0x000CF)]
		'Iuml':                             [rune(0x000CF)]
		'iuml;':                            [rune(0x000EF)]
		'iuml':                             [rune(0x000EF)]
		'Jcirc;':                           [rune(0x00134)]
		'jcirc;':                           [rune(0x00135)]
		'Jcy;':                             [rune(0x00419)]
		'jcy;':                             [rune(0x00439)]
		'Jfr;':                             [rune(0x1D50D)]
		'jfr;':                             [rune(0x1D527)]
		'jmath;':                           [rune(0x00237)]
		'Jopf;':                            [rune(0x1D541)]
		'jopf;':                            [rune(0x1D55B)]
		'Jscr;':                            [rune(0x1D4A5)]
		'jscr;':                            [rune(0x1D4BF)]
		'Jsercy;':                          [rune(0x00408)]
		'jsercy;':                          [rune(0x00458)]
		'Jukcy;':                           [rune(0x00404)]
		'jukcy;':                           [rune(0x00454)]
		'Kappa;':                           [rune(0x0039A)]
		'kappa;':                           [rune(0x003BA)]
		'kappav;':                          [rune(0x003F0)]
		'Kcedil;':                          [rune(0x00136)]
		'kcedil;':                          [rune(0x00137)]
		'Kcy;':                             [rune(0x0041A)]
		'kcy;':                             [rune(0x0043A)]
		'Kfr;':                             [rune(0x1D50E)]
		'kfr;':                             [rune(0x1D528)]
		'kgreen;':                          [rune(0x00138)]
		'KHcy;':                            [rune(0x00425)]
		'khcy;':                            [rune(0x00445)]
		'KJcy;':                            [rune(0x0040C)]
		'kjcy;':                            [rune(0x0045C)]
		'Kopf;':                            [rune(0x1D542)]
		'kopf;':                            [rune(0x1D55C)]
		'Kscr;':                            [rune(0x1D4A6)]
		'kscr;':                            [rune(0x1D4C0)]
		'lAarr;':                           [rune(0x021DA)]
		'Lacute;':                          [rune(0x00139)]
		'lacute;':                          [rune(0x0013A)]
		'laemptyv;':                        [rune(0x029B4)]
		'lagran;':                          [rune(0x02112)]
		'Lambda;':                          [rune(0x0039B)]
		'lambda;':                          [rune(0x003BB)]
		'Lang;':                            [rune(0x027EA)]
		'lang;':                            [rune(0x027E8)]
		'langd;':                           [rune(0x02991)]
		'langle;':                          [rune(0x027E8)]
		'lap;':                             [rune(0x02A85)]
		'Laplacetrf;':                      [rune(0x02112)]
		'laquo;':                           [rune(0x000AB)]
		'laquo':                            [rune(0x000AB)]
		'Larr;':                            [rune(0x0219E)]
		'lArr;':                            [rune(0x021D0)]
		'larr;':                            [rune(0x02190)]
		'larrb;':                           [rune(0x021E4)]
		'larrbfs;':                         [rune(0x0291F)]
		'larrfs;':                          [rune(0x0291D)]
		'larrhk;':                          [rune(0x021A9)]
		'larrlp;':                          [rune(0x021AB)]
		'larrpl;':                          [rune(0x02939)]
		'larrsim;':                         [rune(0x02973)]
		'larrtl;':                          [rune(0x021A2)]
		'lat;':                             [rune(0x02AAB)]
		'lAtail;':                          [rune(0x0291B)]
		'latail;':                          [rune(0x02919)]
		'late;':                            [rune(0x02AAD)]
		'lates;':                           [rune(0x02AAD), 0x0FE00]
		'lBarr;':                           [rune(0x0290E)]
		'lbarr;':                           [rune(0x0290C)]
		'lbbrk;':                           [rune(0x02772)]
		'lbrace;':                          [rune(0x0007B)]
		'lbrack;':                          [rune(0x0005B)]
		'lbrke;':                           [rune(0x0298B)]
		'lbrksld;':                         [rune(0x0298F)]
		'lbrkslu;':                         [rune(0x0298D)]
		'Lcaron;':                          [rune(0x0013D)]
		'lcaron;':                          [rune(0x0013E)]
		'Lcedil;':                          [rune(0x0013B)]
		'lcedil;':                          [rune(0x0013C)]
		'lceil;':                           [rune(0x02308)]
		'lcub;':                            [rune(0x0007B)]
		'Lcy;':                             [rune(0x0041B)]
		'lcy;':                             [rune(0x0043B)]
		'ldca;':                            [rune(0x02936)]
		'ldquo;':                           [rune(0x0201C)]
		'ldquor;':                          [rune(0x0201E)]
		'ldrdhar;':                         [rune(0x02967)]
		'ldrushar;':                        [rune(0x0294B)]
		'ldsh;':                            [rune(0x021B2)]
		'lE;':                              [rune(0x02266)]
		'le;':                              [rune(0x02264)]
		'LeftAngleBracket;':                [rune(0x027E8)]
		'LeftArrow;':                       [rune(0x02190)]
		'Leftarrow;':                       [rune(0x021D0)]
		'leftarrow;':                       [rune(0x02190)]
		'LeftArrowBar;':                    [rune(0x021E4)]
		'LeftArrowRightArrow;':             [rune(0x021C6)]
		'leftarrowtail;':                   [rune(0x021A2)]
		'LeftCeiling;':                     [rune(0x02308)]
		'LeftDoubleBracket;':               [rune(0x027E6)]
		'LeftDownTeeVector;':               [rune(0x02961)]
		'LeftDownVector;':                  [rune(0x021C3)]
		'LeftDownVectorBar;':               [rune(0x02959)]
		'LeftFloor;':                       [rune(0x0230A)]
		'leftharpoondown;':                 [rune(0x021BD)]
		'leftharpoonup;':                   [rune(0x021BC)]
		'leftleftarrows;':                  [rune(0x021C7)]
		'LeftRightArrow;':                  [rune(0x02194)]
		'Leftrightarrow;':                  [rune(0x021D4)]
		'leftrightarrow;':                  [rune(0x02194)]
		'leftrightarrows;':                 [rune(0x021C6)]
		'leftrightharpoons;':               [rune(0x021CB)]
		'leftrightsquigarrow;':             [rune(0x021AD)]
		'LeftRightVector;':                 [rune(0x0294E)]
		'LeftTee;':                         [rune(0x022A3)]
		'LeftTeeArrow;':                    [rune(0x021A4)]
		'LeftTeeVector;':                   [rune(0x0295A)]
		'leftthreetimes;':                  [rune(0x022CB)]
		'LeftTriangle;':                    [rune(0x022B2)]
		'LeftTriangleBar;':                 [rune(0x029CF)]
		'LeftTriangleEqual;':               [rune(0x022B4)]
		'LeftUpDownVector;':                [rune(0x02951)]
		'LeftUpTeeVector;':                 [rune(0x02960)]
		'LeftUpVector;':                    [rune(0x021BF)]
		'LeftUpVectorBar;':                 [rune(0x02958)]
		'LeftVector;':                      [rune(0x021BC)]
		'LeftVectorBar;':                   [rune(0x02952)]
		'lEg;':                             [rune(0x02A8B)]
		'leg;':                             [rune(0x022DA)]
		'leq;':                             [rune(0x02264)]
		'leqq;':                            [rune(0x02266)]
		'leqslant;':                        [rune(0x02A7D)]
		'les;':                             [rune(0x02A7D)]
		'lescc;':                           [rune(0x02AA8)]
		'lesdot;':                          [rune(0x02A7F)]
		'lesdoto;':                         [rune(0x02A81)]
		'lesdotor;':                        [rune(0x02A83)]
		'lesg;':                            [rune(0x022DA), 0x0FE00]
		'lesges;':                          [rune(0x02A93)]
		'lessapprox;':                      [rune(0x02A85)]
		'lessdot;':                         [rune(0x022D6)]
		'lesseqgtr;':                       [rune(0x022DA)]
		'lesseqqgtr;':                      [rune(0x02A8B)]
		'LessEqualGreater;':                [rune(0x022DA)]
		'LessFullEqual;':                   [rune(0x02266)]
		'LessGreater;':                     [rune(0x02276)]
		'lessgtr;':                         [rune(0x02276)]
		'LessLess;':                        [rune(0x02AA1)]
		'lesssim;':                         [rune(0x02272)]
		'LessSlantEqual;':                  [rune(0x02A7D)]
		'LessTilde;':                       [rune(0x02272)]
		'lfisht;':                          [rune(0x0297C)]
		'lfloor;':                          [rune(0x0230A)]
		'Lfr;':                             [rune(0x1D50F)]
		'lfr;':                             [rune(0x1D529)]
		'lg;':                              [rune(0x02276)]
		'lgE;':                             [rune(0x02A91)]
		'lHar;':                            [rune(0x02962)]
		'lhard;':                           [rune(0x021BD)]
		'lharu;':                           [rune(0x021BC)]
		'lharul;':                          [rune(0x0296A)]
		'lhblk;':                           [rune(0x02584)]
		'LJcy;':                            [rune(0x00409)]
		'ljcy;':                            [rune(0x00459)]
		'Ll;':                              [rune(0x022D8)]
		'll;':                              [rune(0x0226A)]
		'llarr;':                           [rune(0x021C7)]
		'llcorner;':                        [rune(0x0231E)]
		'Lleftarrow;':                      [rune(0x021DA)]
		'llhard;':                          [rune(0x0296B)]
		'lltri;':                           [rune(0x025FA)]
		'Lmidot;':                          [rune(0x0013F)]
		'lmidot;':                          [rune(0x00140)]
		'lmoust;':                          [rune(0x023B0)]
		'lmoustache;':                      [rune(0x023B0)]
		'lnap;':                            [rune(0x02A89)]
		'lnapprox;':                        [rune(0x02A89)]
		'lnE;':                             [rune(0x02268)]
		'lne;':                             [rune(0x02A87)]
		'lneq;':                            [rune(0x02A87)]
		'lneqq;':                           [rune(0x02268)]
		'lnsim;':                           [rune(0x022E6)]
		'loang;':                           [rune(0x027EC)]
		'loarr;':                           [rune(0x021FD)]
		'lobrk;':                           [rune(0x027E6)]
		'LongLeftArrow;':                   [rune(0x027F5)]
		'Longleftarrow;':                   [rune(0x027F8)]
		'longleftarrow;':                   [rune(0x027F5)]
		'LongLeftRightArrow;':              [rune(0x027F7)]
		'Longleftrightarrow;':              [rune(0x027FA)]
		'longleftrightarrow;':              [rune(0x027F7)]
		'longmapsto;':                      [rune(0x027FC)]
		'LongRightArrow;':                  [rune(0x027F6)]
		'Longrightarrow;':                  [rune(0x027F9)]
		'longrightarrow;':                  [rune(0x027F6)]
		'looparrowleft;':                   [rune(0x021AB)]
		'looparrowright;':                  [rune(0x021AC)]
		'lopar;':                           [rune(0x02985)]
		'Lopf;':                            [rune(0x1D543)]
		'lopf;':                            [rune(0x1D55D)]
		'loplus;':                          [rune(0x02A2D)]
		'lotimes;':                         [rune(0x02A34)]
		'lowast;':                          [rune(0x02217)]
		'lowbar;':                          [rune(0x0005F)]
		'LowerLeftArrow;':                  [rune(0x02199)]
		'LowerRightArrow;':                 [rune(0x02198)]
		'loz;':                             [rune(0x025CA)]
		'lozenge;':                         [rune(0x025CA)]
		'lozf;':                            [rune(0x029EB)]
		'lpar;':                            [rune(0x00028)]
		'lparlt;':                          [rune(0x02993)]
		'lrarr;':                           [rune(0x021C6)]
		'lrcorner;':                        [rune(0x0231F)]
		'lrhar;':                           [rune(0x021CB)]
		'lrhard;':                          [rune(0x0296D)]
		'lrm;':                             [rune(0x0200E)]
		'lrtri;':                           [rune(0x022BF)]
		'lsaquo;':                          [rune(0x02039)]
		'Lscr;':                            [rune(0x02112)]
		'lscr;':                            [rune(0x1D4C1)]
		'Lsh;':                             [rune(0x021B0)]
		'lsh;':                             [rune(0x021B0)]
		'lsim;':                            [rune(0x02272)]
		'lsime;':                           [rune(0x02A8D)]
		'lsimg;':                           [rune(0x02A8F)]
		'lsqb;':                            [rune(0x0005B)]
		'lsquo;':                           [rune(0x02018)]
		'lsquor;':                          [rune(0x0201A)]
		'Lstrok;':                          [rune(0x00141)]
		'lstrok;':                          [rune(0x00142)]
		'LT;':                              [rune(0x0003C)]
		'LT':                               [rune(0x0003C)]
		'Lt;':                              [rune(0x0226A)]
		'lt;':                              [rune(0x0003C)]
		'lt':                               [rune(0x0003C)]
		'ltcc;':                            [rune(0x02AA6)]
		'ltcir;':                           [rune(0x02A79)]
		'ltdot;':                           [rune(0x022D6)]
		'lthree;':                          [rune(0x022CB)]
		'ltimes;':                          [rune(0x022C9)]
		'ltlarr;':                          [rune(0x02976)]
		'ltquest;':                         [rune(0x02A7B)]
		'ltri;':                            [rune(0x025C3)]
		'ltrie;':                           [rune(0x022B4)]
		'ltrif;':                           [rune(0x025C2)]
		'ltrPar;':                          [rune(0x02996)]
		'lurdshar;':                        [rune(0x0294A)]
		'luruhar;':                         [rune(0x02966)]
		'lvertneqq;':                       [rune(0x02268), 0x0FE00]
		'lvnE;':                            [rune(0x02268), 0x0FE00]
		'macr;':                            [rune(0x000AF)]
		'macr':                             [rune(0x000AF)]
		'male;':                            [rune(0x02642)]
		'malt;':                            [rune(0x02720)]
		'maltese;':                         [rune(0x02720)]
		'Map;':                             [rune(0x02905)]
		'map;':                             [rune(0x021A6)]
		'mapsto;':                          [rune(0x021A6)]
		'mapstodown;':                      [rune(0x021A7)]
		'mapstoleft;':                      [rune(0x021A4)]
		'mapstoup;':                        [rune(0x021A5)]
		'marker;':                          [rune(0x025AE)]
		'mcomma;':                          [rune(0x02A29)]
		'Mcy;':                             [rune(0x0041C)]
		'mcy;':                             [rune(0x0043C)]
		'mdash;':                           [rune(0x02014)]
		'mDDot;':                           [rune(0x0223A)]
		'measuredangle;':                   [rune(0x02221)]
		'MediumSpace;':                     [rune(0x0205F)]
		'Mellintrf;':                       [rune(0x02133)]
		'Mfr;':                             [rune(0x1D510)]
		'mfr;':                             [rune(0x1D52A)]
		'mho;':                             [rune(0x02127)]
		'micro;':                           [rune(0x000B5)]
		'micro':                            [rune(0x000B5)]
		'mid;':                             [rune(0x02223)]
		'midast;':                          [rune(0x0002A)]
		'midcir;':                          [rune(0x02AF0)]
		'middot;':                          [rune(0x000B7)]
		'middot':                           [rune(0x000B7)]
		'minus;':                           [rune(0x02212)]
		'minusb;':                          [rune(0x0229F)]
		'minusd;':                          [rune(0x02238)]
		'minusdu;':                         [rune(0x02A2A)]
		'MinusPlus;':                       [rune(0x02213)]
		'mlcp;':                            [rune(0x02ADB)]
		'mldr;':                            [rune(0x02026)]
		'mnplus;':                          [rune(0x02213)]
		'models;':                          [rune(0x022A7)]
		'Mopf;':                            [rune(0x1D544)]
		'mopf;':                            [rune(0x1D55E)]
		'mp;':                              [rune(0x02213)]
		'Mscr;':                            [rune(0x02133)]
		'mscr;':                            [rune(0x1D4C2)]
		'mstpos;':                          [rune(0x0223E)]
		'Mu;':                              [rune(0x0039C)]
		'mu;':                              [rune(0x003BC)]
		'multimap;':                        [rune(0x022B8)]
		'mumap;':                           [rune(0x022B8)]
		'nabla;':                           [rune(0x02207)]
		'Nacute;':                          [rune(0x00143)]
		'nacute;':                          [rune(0x00144)]
		'nang;':                            [rune(0x02220), 0x020D2]
		'nap;':                             [rune(0x02249)]
		'napE;':                            [rune(0x02A70), 0x00338]
		'napid;':                           [rune(0x0224B), 0x00338]
		'napos;':                           [rune(0x00149)]
		'napprox;':                         [rune(0x02249)]
		'natur;':                           [rune(0x0266E)]
		'natural;':                         [rune(0x0266E)]
		'naturals;':                        [rune(0x02115)]
		'nbsp;':                            [rune(0x000A0)]
		'nbsp':                             [rune(0x000A0)]
		'nbump;':                           [rune(0x0224E), 0x00338]
		'nbumpe;':                          [rune(0x0224F), 0x00338]
		'ncap;':                            [rune(0x02A43)]
		'Ncaron;':                          [rune(0x00147)]
		'ncaron;':                          [rune(0x00148)]
		'Ncedil;':                          [rune(0x00145)]
		'ncedil;':                          [rune(0x00146)]
		'ncong;':                           [rune(0x02247)]
		'ncongdot;':                        [rune(0x02A6D), 0x00338]
		'ncup;':                            [rune(0x02A42)]
		'Ncy;':                             [rune(0x0041D)]
		'ncy;':                             [rune(0x0043D)]
		'ndash;':                           [rune(0x02013)]
		'ne;':                              [rune(0x02260)]
		'nearhk;':                          [rune(0x02924)]
		'neArr;':                           [rune(0x021D7)]
		'nearr;':                           [rune(0x02197)]
		'nearrow;':                         [rune(0x02197)]
		'nedot;':                           [rune(0x02250), 0x00338]
		'NegativeMediumSpace;':             [rune(0x0200B)]
		'NegativeThickSpace;':              [rune(0x0200B)]
		'NegativeThinSpace;':               [rune(0x0200B)]
		'NegativeVeryThinSpace;':           [rune(0x0200B)]
		'nequiv;':                          [rune(0x02262)]
		'nesear;':                          [rune(0x02928)]
		'nesim;':                           [rune(0x02242), 0x00338]
		'NestedGreaterGreater;':            [rune(0x0226B)]
		'NestedLessLess;':                  [rune(0x0226A)]
		'NewLine;':                         [rune(0x0000A)]
		'nexist;':                          [rune(0x02204)]
		'nexists;':                         [rune(0x02204)]
		'Nfr;':                             [rune(0x1D511)]
		'nfr;':                             [rune(0x1D52B)]
		'ngE;':                             [rune(0x02267), 0x00338]
		'nge;':                             [rune(0x02271)]
		'ngeq;':                            [rune(0x02271)]
		'ngeqq;':                           [rune(0x02267), 0x00338]
		'ngeqslant;':                       [rune(0x02A7E), 0x00338]
		'nges;':                            [rune(0x02A7E), 0x00338]
		'nGg;':                             [rune(0x022D9), 0x00338]
		'ngsim;':                           [rune(0x02275)]
		'nGt;':                             [rune(0x0226B), 0x020D2]
		'ngt;':                             [rune(0x0226F)]
		'ngtr;':                            [rune(0x0226F)]
		'nGtv;':                            [rune(0x0226B), 0x00338]
		'nhArr;':                           [rune(0x021CE)]
		'nharr;':                           [rune(0x021AE)]
		'nhpar;':                           [rune(0x02AF2)]
		'ni;':                              [rune(0x0220B)]
		'nis;':                             [rune(0x022FC)]
		'nisd;':                            [rune(0x022FA)]
		'niv;':                             [rune(0x0220B)]
		'NJcy;':                            [rune(0x0040A)]
		'njcy;':                            [rune(0x0045A)]
		'nlArr;':                           [rune(0x021CD)]
		'nlarr;':                           [rune(0x0219A)]
		'nldr;':                            [rune(0x02025)]
		'nlE;':                             [rune(0x02266), 0x00338]
		'nle;':                             [rune(0x02270)]
		'nLeftarrow;':                      [rune(0x021CD)]
		'nleftarrow;':                      [rune(0x0219A)]
		'nLeftrightarrow;':                 [rune(0x021CE)]
		'nleftrightarrow;':                 [rune(0x021AE)]
		'nleq;':                            [rune(0x02270)]
		'nleqq;':                           [rune(0x02266), 0x00338]
		'nleqslant;':                       [rune(0x02A7D), 0x00338]
		'nles;':                            [rune(0x02A7D), 0x00338]
		'nless;':                           [rune(0x0226E)]
		'nLl;':                             [rune(0x022D8), 0x00338]
		'nlsim;':                           [rune(0x02274)]
		'nLt;':                             [rune(0x0226A), 0x020D2]
		'nlt;':                             [rune(0x0226E)]
		'nltri;':                           [rune(0x022EA)]
		'nltrie;':                          [rune(0x022EC)]
		'nLtv;':                            [rune(0x0226A), 0x00338]
		'nmid;':                            [rune(0x02224)]
		'NoBreak;':                         [rune(0x02060)]
		'NonBreakingSpace;':                [rune(0x000A0)]
		'Nopf;':                            [rune(0x02115)]
		'nopf;':                            [rune(0x1D55F)]
		'Not;':                             [rune(0x02AEC)]
		'not;':                             [rune(0x000AC)]
		'not':                              [rune(0x000AC)]
		'NotCongruent;':                    [rune(0x02262)]
		'NotCupCap;':                       [rune(0x0226D)]
		'NotDoubleVerticalBar;':            [rune(0x02226)]
		'NotElement;':                      [rune(0x02209)]
		'NotEqual;':                        [rune(0x02260)]
		'NotEqualTilde;':                   [rune(0x02242), 0x00338]
		'NotExists;':                       [rune(0x02204)]
		'NotGreater;':                      [rune(0x0226F)]
		'NotGreaterEqual;':                 [rune(0x02271)]
		'NotGreaterFullEqual;':             [rune(0x02267), 0x00338]
		'NotGreaterGreater;':               [rune(0x0226B), 0x00338]
		'NotGreaterLess;':                  [rune(0x02279)]
		'NotGreaterSlantEqual;':            [rune(0x02A7E), 0x00338]
		'NotGreaterTilde;':                 [rune(0x02275)]
		'NotHumpDownHump;':                 [rune(0x0224E), 0x00338]
		'NotHumpEqual;':                    [rune(0x0224F), 0x00338]
		'notin;':                           [rune(0x02209)]
		'notindot;':                        [rune(0x022F5), 0x00338]
		'notinE;':                          [rune(0x022F9), 0x00338]
		'notinva;':                         [rune(0x02209)]
		'notinvb;':                         [rune(0x022F7)]
		'notinvc;':                         [rune(0x022F6)]
		'NotLeftTriangle;':                 [rune(0x022EA)]
		'NotLeftTriangleBar;':              [rune(0x029CF), 0x00338]
		'NotLeftTriangleEqual;':            [rune(0x022EC)]
		'NotLess;':                         [rune(0x0226E)]
		'NotLessEqual;':                    [rune(0x02270)]
		'NotLessGreater;':                  [rune(0x02278)]
		'NotLessLess;':                     [rune(0x0226A), 0x00338]
		'NotLessSlantEqual;':               [rune(0x02A7D), 0x00338]
		'NotLessTilde;':                    [rune(0x02274)]
		'NotNestedGreaterGreater;':         [rune(0x02AA2), 0x00338]
		'NotNestedLessLess;':               [rune(0x02AA1), 0x00338]
		'notni;':                           [rune(0x0220C)]
		'notniva;':                         [rune(0x0220C)]
		'notnivb;':                         [rune(0x022FE)]
		'notnivc;':                         [rune(0x022FD)]
		'NotPrecedes;':                     [rune(0x02280)]
		'NotPrecedesEqual;':                [rune(0x02AAF), 0x00338]
		'NotPrecedesSlantEqual;':           [rune(0x022E0)]
		'NotReverseElement;':               [rune(0x0220C)]
		'NotRightTriangle;':                [rune(0x022EB)]
		'NotRightTriangleBar;':             [rune(0x029D0), 0x00338]
		'NotRightTriangleEqual;':           [rune(0x022ED)]
		'NotSquareSubset;':                 [rune(0x0228F), 0x00338]
		'NotSquareSubsetEqual;':            [rune(0x022E2)]
		'NotSquareSuperset;':               [rune(0x02290), 0x00338]
		'NotSquareSupersetEqual;':          [rune(0x022E3)]
		'NotSubset;':                       [rune(0x02282), 0x020D2]
		'NotSubsetEqual;':                  [rune(0x02288)]
		'NotSucceeds;':                     [rune(0x02281)]
		'NotSucceedsEqual;':                [rune(0x02AB0), 0x00338]
		'NotSucceedsSlantEqual;':           [rune(0x022E1)]
		'NotSucceedsTilde;':                [rune(0x0227F), 0x00338]
		'NotSuperset;':                     [rune(0x02283), 0x020D2]
		'NotSupersetEqual;':                [rune(0x02289)]
		'NotTilde;':                        [rune(0x02241)]
		'NotTildeEqual;':                   [rune(0x02244)]
		'NotTildeFullEqual;':               [rune(0x02247)]
		'NotTildeTilde;':                   [rune(0x02249)]
		'NotVerticalBar;':                  [rune(0x02224)]
		'npar;':                            [rune(0x02226)]
		'nparallel;':                       [rune(0x02226)]
		'nparsl;':                          [rune(0x02AFD), 0x020E5]
		'npart;':                           [rune(0x02202), 0x00338]
		'npolint;':                         [rune(0x02A14)]
		'npr;':                             [rune(0x02280)]
		'nprcue;':                          [rune(0x022E0)]
		'npre;':                            [rune(0x02AAF), 0x00338]
		'nprec;':                           [rune(0x02280)]
		'npreceq;':                         [rune(0x02AAF), 0x00338]
		'nrArr;':                           [rune(0x021CF)]
		'nrarr;':                           [rune(0x0219B)]
		'nrarrc;':                          [rune(0x02933), 0x00338]
		'nrarrw;':                          [rune(0x0219D), 0x00338]
		'nRightarrow;':                     [rune(0x021CF)]
		'nrightarrow;':                     [rune(0x0219B)]
		'nrtri;':                           [rune(0x022EB)]
		'nrtrie;':                          [rune(0x022ED)]
		'nsc;':                             [rune(0x02281)]
		'nsccue;':                          [rune(0x022E1)]
		'nsce;':                            [rune(0x02AB0), 0x00338]
		'Nscr;':                            [rune(0x1D4A9)]
		'nscr;':                            [rune(0x1D4C3)]
		'nshortmid;':                       [rune(0x02224)]
		'nshortparallel;':                  [rune(0x02226)]
		'nsim;':                            [rune(0x02241)]
		'nsime;':                           [rune(0x02244)]
		'nsimeq;':                          [rune(0x02244)]
		'nsmid;':                           [rune(0x02224)]
		'nspar;':                           [rune(0x02226)]
		'nsqsube;':                         [rune(0x022E2)]
		'nsqsupe;':                         [rune(0x022E3)]
		'nsub;':                            [rune(0x02284)]
		'nsubE;':                           [rune(0x02AC5), 0x00338]
		'nsube;':                           [rune(0x02288)]
		'nsubset;':                         [rune(0x02282), 0x020D2]
		'nsubseteq;':                       [rune(0x02288)]
		'nsubseteqq;':                      [rune(0x02AC5), 0x00338]
		'nsucc;':                           [rune(0x02281)]
		'nsucceq;':                         [rune(0x02AB0), 0x00338]
		'nsup;':                            [rune(0x02285)]
		'nsupE;':                           [rune(0x02AC6), 0x00338]
		'nsupe;':                           [rune(0x02289)]
		'nsupset;':                         [rune(0x02283), 0x020D2]
		'nsupseteq;':                       [rune(0x02289)]
		'nsupseteqq;':                      [rune(0x02AC6), 0x00338]
		'ntgl;':                            [rune(0x02279)]
		'Ntilde;':                          [rune(0x000D1)]
		'Ntilde':                           [rune(0x000D1)]
		'ntilde;':                          [rune(0x000F1)]
		'ntilde':                           [rune(0x000F1)]
		'ntlg;':                            [rune(0x02278)]
		'ntriangleleft;':                   [rune(0x022EA)]
		'ntrianglelefteq;':                 [rune(0x022EC)]
		'ntriangleright;':                  [rune(0x022EB)]
		'ntrianglerighteq;':                [rune(0x022ED)]
		'Nu;':                              [rune(0x0039D)]
		'nu;':                              [rune(0x003BD)]
		'num;':                             [rune(0x00023)]
		'numero;':                          [rune(0x02116)]
		'numsp;':                           [rune(0x02007)]
		'nvap;':                            [rune(0x0224D), 0x020D2]
		'nVDash;':                          [rune(0x022AF)]
		'nVdash;':                          [rune(0x022AE)]
		'nvDash;':                          [rune(0x022AD)]
		'nvdash;':                          [rune(0x022AC)]
		'nvge;':                            [rune(0x02265), 0x020D2]
		'nvgt;':                            [rune(0x0003E), 0x020D2]
		'nvHarr;':                          [rune(0x02904)]
		'nvinfin;':                         [rune(0x029DE)]
		'nvlArr;':                          [rune(0x02902)]
		'nvle;':                            [rune(0x02264), 0x020D2]
		'nvlt;':                            [rune(0x0003C), 0x020D2]
		'nvltrie;':                         [rune(0x022B4), 0x020D2]
		'nvrArr;':                          [rune(0x02903)]
		'nvrtrie;':                         [rune(0x022B5), 0x020D2]
		'nvsim;':                           [rune(0x0223C), 0x020D2]
		'nwarhk;':                          [rune(0x02923)]
		'nwArr;':                           [rune(0x021D6)]
		'nwarr;':                           [rune(0x02196)]
		'nwarrow;':                         [rune(0x02196)]
		'nwnear;':                          [rune(0x02927)]
		'Oacute;':                          [rune(0x000D3)]
		'Oacute':                           [rune(0x000D3)]
		'oacute;':                          [rune(0x000F3)]
		'oacute':                           [rune(0x000F3)]
		'oast;':                            [rune(0x0229B)]
		'ocir;':                            [rune(0x0229A)]
		'Ocirc;':                           [rune(0x000D4)]
		'Ocirc':                            [rune(0x000D4)]
		'ocirc;':                           [rune(0x000F4)]
		'ocirc':                            [rune(0x000F4)]
		'Ocy;':                             [rune(0x0041E)]
		'ocy;':                             [rune(0x0043E)]
		'odash;':                           [rune(0x0229D)]
		'Odblac;':                          [rune(0x00150)]
		'odblac;':                          [rune(0x00151)]
		'odiv;':                            [rune(0x02A38)]
		'odot;':                            [rune(0x02299)]
		'odsold;':                          [rune(0x029BC)]
		'OElig;':                           [rune(0x00152)]
		'oelig;':                           [rune(0x00153)]
		'ofcir;':                           [rune(0x029BF)]
		'Ofr;':                             [rune(0x1D512)]
		'ofr;':                             [rune(0x1D52C)]
		'ogon;':                            [rune(0x002DB)]
		'Ograve;':                          [rune(0x000D2)]
		'Ograve':                           [rune(0x000D2)]
		'ograve;':                          [rune(0x000F2)]
		'ograve':                           [rune(0x000F2)]
		'ogt;':                             [rune(0x029C1)]
		'ohbar;':                           [rune(0x029B5)]
		'ohm;':                             [rune(0x003A9)]
		'oint;':                            [rune(0x0222E)]
		'olarr;':                           [rune(0x021BA)]
		'olcir;':                           [rune(0x029BE)]
		'olcross;':                         [rune(0x029BB)]
		'oline;':                           [rune(0x0203E)]
		'olt;':                             [rune(0x029C0)]
		'Omacr;':                           [rune(0x0014C)]
		'omacr;':                           [rune(0x0014D)]
		'Omega;':                           [rune(0x003A9)]
		'omega;':                           [rune(0x003C9)]
		'Omicron;':                         [rune(0x0039F)]
		'omicron;':                         [rune(0x003BF)]
		'omid;':                            [rune(0x029B6)]
		'ominus;':                          [rune(0x02296)]
		'Oopf;':                            [rune(0x1D546)]
		'oopf;':                            [rune(0x1D560)]
		'opar;':                            [rune(0x029B7)]
		'OpenCurlyDoubleQuote;':            [rune(0x0201C)]
		'OpenCurlyQuote;':                  [rune(0x02018)]
		'operp;':                           [rune(0x029B9)]
		'oplus;':                           [rune(0x02295)]
		'Or;':                              [rune(0x02A54)]
		'or;':                              [rune(0x02228)]
		'orarr;':                           [rune(0x021BB)]
		'ord;':                             [rune(0x02A5D)]
		'order;':                           [rune(0x02134)]
		'orderof;':                         [rune(0x02134)]
		'ordf;':                            [rune(0x000AA)]
		'ordf':                             [rune(0x000AA)]
		'ordm;':                            [rune(0x000BA)]
		'ordm':                             [rune(0x000BA)]
		'origof;':                          [rune(0x022B6)]
		'oror;':                            [rune(0x02A56)]
		'orslope;':                         [rune(0x02A57)]
		'orv;':                             [rune(0x02A5B)]
		'oS;':                              [rune(0x024C8)]
		'Oscr;':                            [rune(0x1D4AA)]
		'oscr;':                            [rune(0x02134)]
		'Oslash;':                          [rune(0x000D8)]
		'Oslash':                           [rune(0x000D8)]
		'oslash;':                          [rune(0x000F8)]
		'oslash':                           [rune(0x000F8)]
		'osol;':                            [rune(0x02298)]
		'Otilde;':                          [rune(0x000D5)]
		'Otilde':                           [rune(0x000D5)]
		'otilde;':                          [rune(0x000F5)]
		'otilde':                           [rune(0x000F5)]
		'Otimes;':                          [rune(0x02A37)]
		'otimes;':                          [rune(0x02297)]
		'otimesas;':                        [rune(0x02A36)]
		'Ouml;':                            [rune(0x000D6)]
		'Ouml':                             [rune(0x000D6)]
		'ouml;':                            [rune(0x000F6)]
		'ouml':                             [rune(0x000F6)]
		'ovbar;':                           [rune(0x0233D)]
		'OverBar;':                         [rune(0x0203E)]
		'OverBrace;':                       [rune(0x023DE)]
		'OverBracket;':                     [rune(0x023B4)]
		'OverParenthesis;':                 [rune(0x023DC)]
		'par;':                             [rune(0x02225)]
		'para;':                            [rune(0x000B6)]
		'para':                             [rune(0x000B6)]
		'parallel;':                        [rune(0x02225)]
		'parsim;':                          [rune(0x02AF3)]
		'parsl;':                           [rune(0x02AFD)]
		'part;':                            [rune(0x02202)]
		'PartialD;':                        [rune(0x02202)]
		'Pcy;':                             [rune(0x0041F)]
		'pcy;':                             [rune(0x0043F)]
		'percnt;':                          [rune(0x00025)]
		'period;':                          [rune(0x0002E)]
		'permil;':                          [rune(0x02030)]
		'perp;':                            [rune(0x022A5)]
		'pertenk;':                         [rune(0x02031)]
		'Pfr;':                             [rune(0x1D513)]
		'pfr;':                             [rune(0x1D52D)]
		'Phi;':                             [rune(0x003A6)]
		'phi;':                             [rune(0x003C6)]
		'phiv;':                            [rune(0x003D5)]
		'phmmat;':                          [rune(0x02133)]
		'phone;':                           [rune(0x0260E)]
		'Pi;':                              [rune(0x003A0)]
		'pi;':                              [rune(0x003C0)]
		'pitchfork;':                       [rune(0x022D4)]
		'piv;':                             [rune(0x003D6)]
		'planck;':                          [rune(0x0210F)]
		'planckh;':                         [rune(0x0210E)]
		'plankv;':                          [rune(0x0210F)]
		'plus;':                            [rune(0x0002B)]
		'plusacir;':                        [rune(0x02A23)]
		'plusb;':                           [rune(0x0229E)]
		'pluscir;':                         [rune(0x02A22)]
		'plusdo;':                          [rune(0x02214)]
		'plusdu;':                          [rune(0x02A25)]
		'pluse;':                           [rune(0x02A72)]
		'PlusMinus;':                       [rune(0x000B1)]
		'plusmn;':                          [rune(0x000B1)]
		'plusmn':                           [rune(0x000B1)]
		'plussim;':                         [rune(0x02A26)]
		'plustwo;':                         [rune(0x02A27)]
		'pm;':                              [rune(0x000B1)]
		'Poincareplane;':                   [rune(0x0210C)]
		'pointint;':                        [rune(0x02A15)]
		'Popf;':                            [rune(0x02119)]
		'popf;':                            [rune(0x1D561)]
		'pound;':                           [rune(0x000A3)]
		'pound':                            [rune(0x000A3)]
		'Pr;':                              [rune(0x02ABB)]
		'pr;':                              [rune(0x0227A)]
		'prap;':                            [rune(0x02AB7)]
		'prcue;':                           [rune(0x0227C)]
		'prE;':                             [rune(0x02AB3)]
		'pre;':                             [rune(0x02AAF)]
		'prec;':                            [rune(0x0227A)]
		'precapprox;':                      [rune(0x02AB7)]
		'preccurlyeq;':                     [rune(0x0227C)]
		'Precedes;':                        [rune(0x0227A)]
		'PrecedesEqual;':                   [rune(0x02AAF)]
		'PrecedesSlantEqual;':              [rune(0x0227C)]
		'PrecedesTilde;':                   [rune(0x0227E)]
		'preceq;':                          [rune(0x02AAF)]
		'precnapprox;':                     [rune(0x02AB9)]
		'precneqq;':                        [rune(0x02AB5)]
		'precnsim;':                        [rune(0x022E8)]
		'precsim;':                         [rune(0x0227E)]
		'Prime;':                           [rune(0x02033)]
		'prime;':                           [rune(0x02032)]
		'primes;':                          [rune(0x02119)]
		'prnap;':                           [rune(0x02AB9)]
		'prnE;':                            [rune(0x02AB5)]
		'prnsim;':                          [rune(0x022E8)]
		'prod;':                            [rune(0x0220F)]
		'Product;':                         [rune(0x0220F)]
		'profalar;':                        [rune(0x0232E)]
		'profline;':                        [rune(0x02312)]
		'profsurf;':                        [rune(0x02313)]
		'prop;':                            [rune(0x0221D)]
		'Proportion;':                      [rune(0x02237)]
		'Proportional;':                    [rune(0x0221D)]
		'propto;':                          [rune(0x0221D)]
		'prsim;':                           [rune(0x0227E)]
		'prurel;':                          [rune(0x022B0)]
		'Pscr;':                            [rune(0x1D4AB)]
		'pscr;':                            [rune(0x1D4C5)]
		'Psi;':                             [rune(0x003A8)]
		'psi;':                             [rune(0x003C8)]
		'puncsp;':                          [rune(0x02008)]
		'Qfr;':                             [rune(0x1D514)]
		'qfr;':                             [rune(0x1D52E)]
		'qint;':                            [rune(0x02A0C)]
		'Qopf;':                            [rune(0x0211A)]
		'qopf;':                            [rune(0x1D562)]
		'qprime;':                          [rune(0x02057)]
		'Qscr;':                            [rune(0x1D4AC)]
		'qscr;':                            [rune(0x1D4C6)]
		'quaternions;':                     [rune(0x0210D)]
		'quatint;':                         [rune(0x02A16)]
		'quest;':                           [rune(0x0003F)]
		'questeq;':                         [rune(0x0225F)]
		'QUOT;':                            [rune(0x00022)]
		'QUOT':                             [rune(0x00022)]
		'quot;':                            [rune(0x00022)]
		'quot':                             [rune(0x00022)]
		'rAarr;':                           [rune(0x021DB)]
		'race;':                            [rune(0x0223D), 0x00331]
		'Racute;':                          [rune(0x00154)]
		'racute;':                          [rune(0x00155)]
		'radic;':                           [rune(0x0221A)]
		'raemptyv;':                        [rune(0x029B3)]
		'Rang;':                            [rune(0x027EB)]
		'rang;':                            [rune(0x027E9)]
		'rangd;':                           [rune(0x02992)]
		'range;':                           [rune(0x029A5)]
		'rangle;':                          [rune(0x027E9)]
		'raquo;':                           [rune(0x000BB)]
		'raquo':                            [rune(0x000BB)]
		'Rarr;':                            [rune(0x021A0)]
		'rArr;':                            [rune(0x021D2)]
		'rarr;':                            [rune(0x02192)]
		'rarrap;':                          [rune(0x02975)]
		'rarrb;':                           [rune(0x021E5)]
		'rarrbfs;':                         [rune(0x02920)]
		'rarrc;':                           [rune(0x02933)]
		'rarrfs;':                          [rune(0x0291E)]
		'rarrhk;':                          [rune(0x021AA)]
		'rarrlp;':                          [rune(0x021AC)]
		'rarrpl;':                          [rune(0x02945)]
		'rarrsim;':                         [rune(0x02974)]
		'Rarrtl;':                          [rune(0x02916)]
		'rarrtl;':                          [rune(0x021A3)]
		'rarrw;':                           [rune(0x0219D)]
		'rAtail;':                          [rune(0x0291C)]
		'ratail;':                          [rune(0x0291A)]
		'ratio;':                           [rune(0x02236)]
		'rationals;':                       [rune(0x0211A)]
		'RBarr;':                           [rune(0x02910)]
		'rBarr;':                           [rune(0x0290F)]
		'rbarr;':                           [rune(0x0290D)]
		'rbbrk;':                           [rune(0x02773)]
		'rbrace;':                          [rune(0x0007D)]
		'rbrack;':                          [rune(0x0005D)]
		'rbrke;':                           [rune(0x0298C)]
		'rbrksld;':                         [rune(0x0298E)]
		'rbrkslu;':                         [rune(0x02990)]
		'Rcaron;':                          [rune(0x00158)]
		'rcaron;':                          [rune(0x00159)]
		'Rcedil;':                          [rune(0x00156)]
		'rcedil;':                          [rune(0x00157)]
		'rceil;':                           [rune(0x02309)]
		'rcub;':                            [rune(0x0007D)]
		'Rcy;':                             [rune(0x00420)]
		'rcy;':                             [rune(0x00440)]
		'rdca;':                            [rune(0x02937)]
		'rdldhar;':                         [rune(0x02969)]
		'rdquo;':                           [rune(0x0201D)]
		'rdquor;':                          [rune(0x0201D)]
		'rdsh;':                            [rune(0x021B3)]
		'Re;':                              [rune(0x0211C)]
		'real;':                            [rune(0x0211C)]
		'realine;':                         [rune(0x0211B)]
		'realpart;':                        [rune(0x0211C)]
		'reals;':                           [rune(0x0211D)]
		'rect;':                            [rune(0x025AD)]
		'REG;':                             [rune(0x000AE)]
		'REG':                              [rune(0x000AE)]
		'reg;':                             [rune(0x000AE)]
		'reg':                              [rune(0x000AE)]
		'ReverseElement;':                  [rune(0x0220B)]
		'ReverseEquilibrium;':              [rune(0x021CB)]
		'ReverseUpEquilibrium;':            [rune(0x0296F)]
		'rfisht;':                          [rune(0x0297D)]
		'rfloor;':                          [rune(0x0230B)]
		'Rfr;':                             [rune(0x0211C)]
		'rfr;':                             [rune(0x1D52F)]
		'rHar;':                            [rune(0x02964)]
		'rhard;':                           [rune(0x021C1)]
		'rharu;':                           [rune(0x021C0)]
		'rharul;':                          [rune(0x0296C)]
		'Rho;':                             [rune(0x003A1)]
		'rho;':                             [rune(0x003C1)]
		'rhov;':                            [rune(0x003F1)]
		'RightAngleBracket;':               [rune(0x027E9)]
		'RightArrow;':                      [rune(0x02192)]
		'Rightarrow;':                      [rune(0x021D2)]
		'rightarrow;':                      [rune(0x02192)]
		'RightArrowBar;':                   [rune(0x021E5)]
		'RightArrowLeftArrow;':             [rune(0x021C4)]
		'rightarrowtail;':                  [rune(0x021A3)]
		'RightCeiling;':                    [rune(0x02309)]
		'RightDoubleBracket;':              [rune(0x027E7)]
		'RightDownTeeVector;':              [rune(0x0295D)]
		'RightDownVector;':                 [rune(0x021C2)]
		'RightDownVectorBar;':              [rune(0x02955)]
		'RightFloor;':                      [rune(0x0230B)]
		'rightharpoondown;':                [rune(0x021C1)]
		'rightharpoonup;':                  [rune(0x021C0)]
		'rightleftarrows;':                 [rune(0x021C4)]
		'rightleftharpoons;':               [rune(0x021CC)]
		'rightrightarrows;':                [rune(0x021C9)]
		'rightsquigarrow;':                 [rune(0x0219D)]
		'RightTee;':                        [rune(0x022A2)]
		'RightTeeArrow;':                   [rune(0x021A6)]
		'RightTeeVector;':                  [rune(0x0295B)]
		'rightthreetimes;':                 [rune(0x022CC)]
		'RightTriangle;':                   [rune(0x022B3)]
		'RightTriangleBar;':                [rune(0x029D0)]
		'RightTriangleEqual;':              [rune(0x022B5)]
		'RightUpDownVector;':               [rune(0x0294F)]
		'RightUpTeeVector;':                [rune(0x0295C)]
		'RightUpVector;':                   [rune(0x021BE)]
		'RightUpVectorBar;':                [rune(0x02954)]
		'RightVector;':                     [rune(0x021C0)]
		'RightVectorBar;':                  [rune(0x02953)]
		'ring;':                            [rune(0x002DA)]
		'risingdotseq;':                    [rune(0x02253)]
		'rlarr;':                           [rune(0x021C4)]
		'rlhar;':                           [rune(0x021CC)]
		'rlm;':                             [rune(0x0200F)]
		'rmoust;':                          [rune(0x023B1)]
		'rmoustache;':                      [rune(0x023B1)]
		'rnmid;':                           [rune(0x02AEE)]
		'roang;':                           [rune(0x027ED)]
		'roarr;':                           [rune(0x021FE)]
		'robrk;':                           [rune(0x027E7)]
		'ropar;':                           [rune(0x02986)]
		'Ropf;':                            [rune(0x0211D)]
		'ropf;':                            [rune(0x1D563)]
		'roplus;':                          [rune(0x02A2E)]
		'rotimes;':                         [rune(0x02A35)]
		'RoundImplies;':                    [rune(0x02970)]
		'rpar;':                            [rune(0x00029)]
		'rpargt;':                          [rune(0x02994)]
		'rppolint;':                        [rune(0x02A12)]
		'rrarr;':                           [rune(0x021C9)]
		'Rrightarrow;':                     [rune(0x021DB)]
		'rsaquo;':                          [rune(0x0203A)]
		'Rscr;':                            [rune(0x0211B)]
		'rscr;':                            [rune(0x1D4C7)]
		'Rsh;':                             [rune(0x021B1)]
		'rsh;':                             [rune(0x021B1)]
		'rsqb;':                            [rune(0x0005D)]
		'rsquo;':                           [rune(0x02019)]
		'rsquor;':                          [rune(0x02019)]
		'rthree;':                          [rune(0x022CC)]
		'rtimes;':                          [rune(0x022CA)]
		'rtri;':                            [rune(0x025B9)]
		'rtrie;':                           [rune(0x022B5)]
		'rtrif;':                           [rune(0x025B8)]
		'rtriltri;':                        [rune(0x029CE)]
		'RuleDelayed;':                     [rune(0x029F4)]
		'ruluhar;':                         [rune(0x02968)]
		'rx;':                              [rune(0x0211E)]
		'Sacute;':                          [rune(0x0015A)]
		'sacute;':                          [rune(0x0015B)]
		'sbquo;':                           [rune(0x0201A)]
		'Sc;':                              [rune(0x02ABC)]
		'sc;':                              [rune(0x0227B)]
		'scap;':                            [rune(0x02AB8)]
		'Scaron;':                          [rune(0x00160)]
		'scaron;':                          [rune(0x00161)]
		'sccue;':                           [rune(0x0227D)]
		'scE;':                             [rune(0x02AB4)]
		'sce;':                             [rune(0x02AB0)]
		'Scedil;':                          [rune(0x0015E)]
		'scedil;':                          [rune(0x0015F)]
		'Scirc;':                           [rune(0x0015C)]
		'scirc;':                           [rune(0x0015D)]
		'scnap;':                           [rune(0x02ABA)]
		'scnE;':                            [rune(0x02AB6)]
		'scnsim;':                          [rune(0x022E9)]
		'scpolint;':                        [rune(0x02A13)]
		'scsim;':                           [rune(0x0227F)]
		'Scy;':                             [rune(0x00421)]
		'scy;':                             [rune(0x00441)]
		'sdot;':                            [rune(0x022C5)]
		'sdotb;':                           [rune(0x022A1)]
		'sdote;':                           [rune(0x02A66)]
		'searhk;':                          [rune(0x02925)]
		'seArr;':                           [rune(0x021D8)]
		'searr;':                           [rune(0x02198)]
		'searrow;':                         [rune(0x02198)]
		'sect;':                            [rune(0x000A7)]
		'sect':                             [rune(0x000A7)]
		'semi;':                            [rune(0x0003B)]
		'seswar;':                          [rune(0x02929)]
		'setminus;':                        [rune(0x02216)]
		'setmn;':                           [rune(0x02216)]
		'sext;':                            [rune(0x02736)]
		'Sfr;':                             [rune(0x1D516)]
		'sfr;':                             [rune(0x1D530)]
		'sfrown;':                          [rune(0x02322)]
		'sharp;':                           [rune(0x0266F)]
		'SHCHcy;':                          [rune(0x00429)]
		'shchcy;':                          [rune(0x00449)]
		'SHcy;':                            [rune(0x00428)]
		'shcy;':                            [rune(0x00448)]
		'ShortDownArrow;':                  [rune(0x02193)]
		'ShortLeftArrow;':                  [rune(0x02190)]
		'shortmid;':                        [rune(0x02223)]
		'shortparallel;':                   [rune(0x02225)]
		'ShortRightArrow;':                 [rune(0x02192)]
		'ShortUpArrow;':                    [rune(0x02191)]
		'shy;':                             [rune(0x000AD)]
		'shy':                              [rune(0x000AD)]
		'Sigma;':                           [rune(0x003A3)]
		'sigma;':                           [rune(0x003C3)]
		'sigmaf;':                          [rune(0x003C2)]
		'sigmav;':                          [rune(0x003C2)]
		'sim;':                             [rune(0x0223C)]
		'simdot;':                          [rune(0x02A6A)]
		'sime;':                            [rune(0x02243)]
		'simeq;':                           [rune(0x02243)]
		'simg;':                            [rune(0x02A9E)]
		'simgE;':                           [rune(0x02AA0)]
		'siml;':                            [rune(0x02A9D)]
		'simlE;':                           [rune(0x02A9F)]
		'simne;':                           [rune(0x02246)]
		'simplus;':                         [rune(0x02A24)]
		'simrarr;':                         [rune(0x02972)]
		'slarr;':                           [rune(0x02190)]
		'SmallCircle;':                     [rune(0x02218)]
		'smallsetminus;':                   [rune(0x02216)]
		'smashp;':                          [rune(0x02A33)]
		'smeparsl;':                        [rune(0x029E4)]
		'smid;':                            [rune(0x02223)]
		'smile;':                           [rune(0x02323)]
		'smt;':                             [rune(0x02AAA)]
		'smte;':                            [rune(0x02AAC)]
		'smtes;':                           [rune(0x02AAC), 0x0FE00]
		'SOFTcy;':                          [rune(0x0042C)]
		'softcy;':                          [rune(0x0044C)]
		'sol;':                             [rune(0x0002F)]
		'solb;':                            [rune(0x029C4)]
		'solbar;':                          [rune(0x0233F)]
		'Sopf;':                            [rune(0x1D54A)]
		'sopf;':                            [rune(0x1D564)]
		'spades;':                          [rune(0x02660)]
		'spadesuit;':                       [rune(0x02660)]
		'spar;':                            [rune(0x02225)]
		'sqcap;':                           [rune(0x02293)]
		'sqcaps;':                          [rune(0x02293), 0x0FE00]
		'sqcup;':                           [rune(0x02294)]
		'sqcups;':                          [rune(0x02294), 0x0FE00]
		'Sqrt;':                            [rune(0x0221A)]
		'sqsub;':                           [rune(0x0228F)]
		'sqsube;':                          [rune(0x02291)]
		'sqsubset;':                        [rune(0x0228F)]
		'sqsubseteq;':                      [rune(0x02291)]
		'sqsup;':                           [rune(0x02290)]
		'sqsupe;':                          [rune(0x02292)]
		'sqsupset;':                        [rune(0x02290)]
		'sqsupseteq;':                      [rune(0x02292)]
		'squ;':                             [rune(0x025A1)]
		'Square;':                          [rune(0x025A1)]
		'square;':                          [rune(0x025A1)]
		'SquareIntersection;':              [rune(0x02293)]
		'SquareSubset;':                    [rune(0x0228F)]
		'SquareSubsetEqual;':               [rune(0x02291)]
		'SquareSuperset;':                  [rune(0x02290)]
		'SquareSupersetEqual;':             [rune(0x02292)]
		'SquareUnion;':                     [rune(0x02294)]
		'squarf;':                          [rune(0x025AA)]
		'squf;':                            [rune(0x025AA)]
		'srarr;':                           [rune(0x02192)]
		'Sscr;':                            [rune(0x1D4AE)]
		'sscr;':                            [rune(0x1D4C8)]
		'ssetmn;':                          [rune(0x02216)]
		'ssmile;':                          [rune(0x02323)]
		'sstarf;':                          [rune(0x022C6)]
		'Star;':                            [rune(0x022C6)]
		'star;':                            [rune(0x02606)]
		'starf;':                           [rune(0x02605)]
		'straightepsilon;':                 [rune(0x003F5)]
		'straightphi;':                     [rune(0x003D5)]
		'strns;':                           [rune(0x000AF)]
		'Sub;':                             [rune(0x022D0)]
		'sub;':                             [rune(0x02282)]
		'subdot;':                          [rune(0x02ABD)]
		'subE;':                            [rune(0x02AC5)]
		'sube;':                            [rune(0x02286)]
		'subedot;':                         [rune(0x02AC3)]
		'submult;':                         [rune(0x02AC1)]
		'subnE;':                           [rune(0x02ACB)]
		'subne;':                           [rune(0x0228A)]
		'subplus;':                         [rune(0x02ABF)]
		'subrarr;':                         [rune(0x02979)]
		'Subset;':                          [rune(0x022D0)]
		'subset;':                          [rune(0x02282)]
		'subseteq;':                        [rune(0x02286)]
		'subseteqq;':                       [rune(0x02AC5)]
		'SubsetEqual;':                     [rune(0x02286)]
		'subsetneq;':                       [rune(0x0228A)]
		'subsetneqq;':                      [rune(0x02ACB)]
		'subsim;':                          [rune(0x02AC7)]
		'subsub;':                          [rune(0x02AD5)]
		'subsup;':                          [rune(0x02AD3)]
		'succ;':                            [rune(0x0227B)]
		'succapprox;':                      [rune(0x02AB8)]
		'succcurlyeq;':                     [rune(0x0227D)]
		'Succeeds;':                        [rune(0x0227B)]
		'SucceedsEqual;':                   [rune(0x02AB0)]
		'SucceedsSlantEqual;':              [rune(0x0227D)]
		'SucceedsTilde;':                   [rune(0x0227F)]
		'succeq;':                          [rune(0x02AB0)]
		'succnapprox;':                     [rune(0x02ABA)]
		'succneqq;':                        [rune(0x02AB6)]
		'succnsim;':                        [rune(0x022E9)]
		'succsim;':                         [rune(0x0227F)]
		'SuchThat;':                        [rune(0x0220B)]
		'Sum;':                             [rune(0x02211)]
		'sum;':                             [rune(0x02211)]
		'sung;':                            [rune(0x0266A)]
		'Sup;':                             [rune(0x022D1)]
		'sup;':                             [rune(0x02283)]
		'sup1;':                            [rune(0x000B9)]
		'sup1':                             [rune(0x000B9)]
		'sup2;':                            [rune(0x000B2)]
		'sup2':                             [rune(0x000B2)]
		'sup3;':                            [rune(0x000B3)]
		'sup3':                             [rune(0x000B3)]
		'supdot;':                          [rune(0x02ABE)]
		'supdsub;':                         [rune(0x02AD8)]
		'supE;':                            [rune(0x02AC6)]
		'supe;':                            [rune(0x02287)]
		'supedot;':                         [rune(0x02AC4)]
		'Superset;':                        [rune(0x02283)]
		'SupersetEqual;':                   [rune(0x02287)]
		'suphsol;':                         [rune(0x027C9)]
		'suphsub;':                         [rune(0x02AD7)]
		'suplarr;':                         [rune(0x0297B)]
		'supmult;':                         [rune(0x02AC2)]
		'supnE;':                           [rune(0x02ACC)]
		'supne;':                           [rune(0x0228B)]
		'supplus;':                         [rune(0x02AC0)]
		'Supset;':                          [rune(0x022D1)]
		'supset;':                          [rune(0x02283)]
		'supseteq;':                        [rune(0x02287)]
		'supseteqq;':                       [rune(0x02AC6)]
		'supsetneq;':                       [rune(0x0228B)]
		'supsetneqq;':                      [rune(0x02ACC)]
		'supsim;':                          [rune(0x02AC8)]
		'supsub;':                          [rune(0x02AD4)]
		'supsup;':                          [rune(0x02AD6)]
		'swarhk;':                          [rune(0x02926)]
		'swArr;':                           [rune(0x021D9)]
		'swarr;':                           [rune(0x02199)]
		'swarrow;':                         [rune(0x02199)]
		'swnwar;':                          [rune(0x0292A)]
		'szlig;':                           [rune(0x000DF)]
		'szlig':                            [rune(0x000DF)]
		'Tab;':                             [rune(0x00009)]
		'target;':                          [rune(0x02316)]
		'Tau;':                             [rune(0x003A4)]
		'tau;':                             [rune(0x003C4)]
		'tbrk;':                            [rune(0x023B4)]
		'Tcaron;':                          [rune(0x00164)]
		'tcaron;':                          [rune(0x00165)]
		'Tcedil;':                          [rune(0x00162)]
		'tcedil;':                          [rune(0x00163)]
		'Tcy;':                             [rune(0x00422)]
		'tcy;':                             [rune(0x00442)]
		'tdot;':                            [rune(0x020DB)]
		'telrec;':                          [rune(0x02315)]
		'Tfr;':                             [rune(0x1D517)]
		'tfr;':                             [rune(0x1D531)]
		'there4;':                          [rune(0x02234)]
		'Therefore;':                       [rune(0x02234)]
		'therefore;':                       [rune(0x02234)]
		'Theta;':                           [rune(0x00398)]
		'theta;':                           [rune(0x003B8)]
		'thetasym;':                        [rune(0x003D1)]
		'thetav;':                          [rune(0x003D1)]
		'thickapprox;':                     [rune(0x02248)]
		'thicksim;':                        [rune(0x0223C)]
		'ThickSpace;':                      [rune(0x0205F), 0x0200A]
		'thinsp;':                          [rune(0x02009)]
		'ThinSpace;':                       [rune(0x02009)]
		'thkap;':                           [rune(0x02248)]
		'thksim;':                          [rune(0x0223C)]
		'THORN;':                           [rune(0x000DE)]
		'THORN':                            [rune(0x000DE)]
		'thorn;':                           [rune(0x000FE)]
		'thorn':                            [rune(0x000FE)]
		'Tilde;':                           [rune(0x0223C)]
		'tilde;':                           [rune(0x002DC)]
		'TildeEqual;':                      [rune(0x02243)]
		'TildeFullEqual;':                  [rune(0x02245)]
		'TildeTilde;':                      [rune(0x02248)]
		'times;':                           [rune(0x000D7)]
		'times':                            [rune(0x000D7)]
		'timesb;':                          [rune(0x022A0)]
		'timesbar;':                        [rune(0x02A31)]
		'timesd;':                          [rune(0x02A30)]
		'tint;':                            [rune(0x0222D)]
		'toea;':                            [rune(0x02928)]
		'top;':                             [rune(0x022A4)]
		'topbot;':                          [rune(0x02336)]
		'topcir;':                          [rune(0x02AF1)]
		'Topf;':                            [rune(0x1D54B)]
		'topf;':                            [rune(0x1D565)]
		'topfork;':                         [rune(0x02ADA)]
		'tosa;':                            [rune(0x02929)]
		'tprime;':                          [rune(0x02034)]
		'TRADE;':                           [rune(0x02122)]
		'trade;':                           [rune(0x02122)]
		'triangle;':                        [rune(0x025B5)]
		'triangledown;':                    [rune(0x025BF)]
		'triangleleft;':                    [rune(0x025C3)]
		'trianglelefteq;':                  [rune(0x022B4)]
		'triangleq;':                       [rune(0x0225C)]
		'triangleright;':                   [rune(0x025B9)]
		'trianglerighteq;':                 [rune(0x022B5)]
		'tridot;':                          [rune(0x025EC)]
		'trie;':                            [rune(0x0225C)]
		'triminus;':                        [rune(0x02A3A)]
		'TripleDot;':                       [rune(0x020DB)]
		'triplus;':                         [rune(0x02A39)]
		'trisb;':                           [rune(0x029CD)]
		'tritime;':                         [rune(0x02A3B)]
		'trpezium;':                        [rune(0x023E2)]
		'Tscr;':                            [rune(0x1D4AF)]
		'tscr;':                            [rune(0x1D4C9)]
		'TScy;':                            [rune(0x00426)]
		'tscy;':                            [rune(0x00446)]
		'TSHcy;':                           [rune(0x0040B)]
		'tshcy;':                           [rune(0x0045B)]
		'Tstrok;':                          [rune(0x00166)]
		'tstrok;':                          [rune(0x00167)]
		'twixt;':                           [rune(0x0226C)]
		'twoheadleftarrow;':                [rune(0x0219E)]
		'twoheadrightarrow;':               [rune(0x021A0)]
		'Uacute;':                          [rune(0x000DA)]
		'Uacute':                           [rune(0x000DA)]
		'uacute;':                          [rune(0x000FA)]
		'uacute':                           [rune(0x000FA)]
		'Uarr;':                            [rune(0x0219F)]
		'uArr;':                            [rune(0x021D1)]
		'uarr;':                            [rune(0x02191)]
		'Uarrocir;':                        [rune(0x02949)]
		'Ubrcy;':                           [rune(0x0040E)]
		'ubrcy;':                           [rune(0x0045E)]
		'Ubreve;':                          [rune(0x0016C)]
		'ubreve;':                          [rune(0x0016D)]
		'Ucirc;':                           [rune(0x000DB)]
		'Ucirc':                            [rune(0x000DB)]
		'ucirc;':                           [rune(0x000FB)]
		'ucirc':                            [rune(0x000FB)]
		'Ucy;':                             [rune(0x00423)]
		'ucy;':                             [rune(0x00443)]
		'udarr;':                           [rune(0x021C5)]
		'Udblac;':                          [rune(0x00170)]
		'udblac;':                          [rune(0x00171)]
		'udhar;':                           [rune(0x0296E)]
		'ufisht;':                          [rune(0x0297E)]
		'Ufr;':                             [rune(0x1D518)]
		'ufr;':                             [rune(0x1D532)]
		'Ugrave;':                          [rune(0x000D9)]
		'Ugrave':                           [rune(0x000D9)]
		'ugrave;':                          [rune(0x000F9)]
		'ugrave':                           [rune(0x000F9)]
		'uHar;':                            [rune(0x02963)]
		'uharl;':                           [rune(0x021BF)]
		'uharr;':                           [rune(0x021BE)]
		'uhblk;':                           [rune(0x02580)]
		'ulcorn;':                          [rune(0x0231C)]
		'ulcorner;':                        [rune(0x0231C)]
		'ulcrop;':                          [rune(0x0230F)]
		'ultri;':                           [rune(0x025F8)]
		'Umacr;':                           [rune(0x0016A)]
		'umacr;':                           [rune(0x0016B)]
		'uml;':                             [rune(0x000A8)]
		'uml':                              [rune(0x000A8)]
		'UnderBar;':                        [rune(0x0005F)]
		'UnderBrace;':                      [rune(0x023DF)]
		'UnderBracket;':                    [rune(0x023B5)]
		'UnderParenthesis;':                [rune(0x023DD)]
		'Union;':                           [rune(0x022C3)]
		'UnionPlus;':                       [rune(0x0228E)]
		'Uogon;':                           [rune(0x00172)]
		'uogon;':                           [rune(0x00173)]
		'Uopf;':                            [rune(0x1D54C)]
		'uopf;':                            [rune(0x1D566)]
		'UpArrow;':                         [rune(0x02191)]
		'Uparrow;':                         [rune(0x021D1)]
		'uparrow;':                         [rune(0x02191)]
		'UpArrowBar;':                      [rune(0x02912)]
		'UpArrowDownArrow;':                [rune(0x021C5)]
		'UpDownArrow;':                     [rune(0x02195)]
		'Updownarrow;':                     [rune(0x021D5)]
		'updownarrow;':                     [rune(0x02195)]
		'UpEquilibrium;':                   [rune(0x0296E)]
		'upharpoonleft;':                   [rune(0x021BF)]
		'upharpoonright;':                  [rune(0x021BE)]
		'uplus;':                           [rune(0x0228E)]
		'UpperLeftArrow;':                  [rune(0x02196)]
		'UpperRightArrow;':                 [rune(0x02197)]
		'Upsi;':                            [rune(0x003D2)]
		'upsi;':                            [rune(0x003C5)]
		'upsih;':                           [rune(0x003D2)]
		'Upsilon;':                         [rune(0x003A5)]
		'upsilon;':                         [rune(0x003C5)]
		'UpTee;':                           [rune(0x022A5)]
		'UpTeeArrow;':                      [rune(0x021A5)]
		'upuparrows;':                      [rune(0x021C8)]
		'urcorn;':                          [rune(0x0231D)]
		'urcorner;':                        [rune(0x0231D)]
		'urcrop;':                          [rune(0x0230E)]
		'Uring;':                           [rune(0x0016E)]
		'uring;':                           [rune(0x0016F)]
		'urtri;':                           [rune(0x025F9)]
		'Uscr;':                            [rune(0x1D4B0)]
		'uscr;':                            [rune(0x1D4CA)]
		'utdot;':                           [rune(0x022F0)]
		'Utilde;':                          [rune(0x00168)]
		'utilde;':                          [rune(0x00169)]
		'utri;':                            [rune(0x025B5)]
		'utrif;':                           [rune(0x025B4)]
		'uuarr;':                           [rune(0x021C8)]
		'Uuml;':                            [rune(0x000DC)]
		'Uuml':                             [rune(0x000DC)]
		'uuml;':                            [rune(0x000FC)]
		'uuml':                             [rune(0x000FC)]
		'uwangle;':                         [rune(0x029A7)]
		'vangrt;':                          [rune(0x0299C)]
		'varepsilon;':                      [rune(0x003F5)]
		'varkappa;':                        [rune(0x003F0)]
		'varnothing;':                      [rune(0x02205)]
		'varphi;':                          [rune(0x003D5)]
		'varpi;':                           [rune(0x003D6)]
		'varpropto;':                       [rune(0x0221D)]
		'vArr;':                            [rune(0x021D5)]
		'varr;':                            [rune(0x02195)]
		'varrho;':                          [rune(0x003F1)]
		'varsigma;':                        [rune(0x003C2)]
		'varsubsetneq;':                    [rune(0x0228A), 0x0FE00]
		'varsubsetneqq;':                   [rune(0x02ACB), 0x0FE00]
		'varsupsetneq;':                    [rune(0x0228B), 0x0FE00]
		'varsupsetneqq;':                   [rune(0x02ACC), 0x0FE00]
		'vartheta;':                        [rune(0x003D1)]
		'vartriangleleft;':                 [rune(0x022B2)]
		'vartriangleright;':                [rune(0x022B3)]
		'Vbar;':                            [rune(0x02AEB)]
		'vBar;':                            [rune(0x02AE8)]
		'vBarv;':                           [rune(0x02AE9)]
		'Vcy;':                             [rune(0x00412)]
		'vcy;':                             [rune(0x00432)]
		'VDash;':                           [rune(0x022AB)]
		'Vdash;':                           [rune(0x022A9)]
		'vDash;':                           [rune(0x022A8)]
		'vdash;':                           [rune(0x022A2)]
		'Vdashl;':                          [rune(0x02AE6)]
		'Vee;':                             [rune(0x022C1)]
		'vee;':                             [rune(0x02228)]
		'veebar;':                          [rune(0x022BB)]
		'veeeq;':                           [rune(0x0225A)]
		'vellip;':                          [rune(0x022EE)]
		'Verbar;':                          [rune(0x02016)]
		'verbar;':                          [rune(0x0007C)]
		'Vert;':                            [rune(0x02016)]
		'vert;':                            [rune(0x0007C)]
		'VerticalBar;':                     [rune(0x02223)]
		'VerticalLine;':                    [rune(0x0007C)]
		'VerticalSeparator;':               [rune(0x02758)]
		'VerticalTilde;':                   [rune(0x02240)]
		'VeryThinSpace;':                   [rune(0x0200A)]
		'Vfr;':                             [rune(0x1D519)]
		'vfr;':                             [rune(0x1D533)]
		'vltri;':                           [rune(0x022B2)]
		'vnsub;':                           [rune(0x02282), 0x020D2]
		'vnsup;':                           [rune(0x02283), 0x020D2]
		'Vopf;':                            [rune(0x1D54D)]
		'vopf;':                            [rune(0x1D567)]
		'vprop;':                           [rune(0x0221D)]
		'vrtri;':                           [rune(0x022B3)]
		'Vscr;':                            [rune(0x1D4B1)]
		'vscr;':                            [rune(0x1D4CB)]
		'vsubnE;':                          [rune(0x02ACB), 0x0FE00]
		'vsubne;':                          [rune(0x0228A), 0x0FE00]
		'vsupnE;':                          [rune(0x02ACC), 0x0FE00]
		'vsupne;':                          [rune(0x0228B), 0x0FE00]
		'Vvdash;':                          [rune(0x022AA)]
		'vzigzag;':                         [rune(0x0299A)]
		'Wcirc;':                           [rune(0x00174)]
		'wcirc;':                           [rune(0x00175)]
		'wedbar;':                          [rune(0x02A5F)]
		'Wedge;':                           [rune(0x022C0)]
		'wedge;':                           [rune(0x02227)]
		'wedgeq;':                          [rune(0x02259)]
		'weierp;':                          [rune(0x02118)]
		'Wfr;':                             [rune(0x1D51A)]
		'wfr;':                             [rune(0x1D534)]
		'Wopf;':                            [rune(0x1D54E)]
		'wopf;':                            [rune(0x1D568)]
		'wp;':                              [rune(0x02118)]
		'wr;':                              [rune(0x02240)]
		'wreath;':                          [rune(0x02240)]
		'Wscr;':                            [rune(0x1D4B2)]
		'wscr;':                            [rune(0x1D4CC)]
		'xcap;':                            [rune(0x022C2)]
		'xcirc;':                           [rune(0x025EF)]
		'xcup;':                            [rune(0x022C3)]
		'xdtri;':                           [rune(0x025BD)]
		'Xfr;':                             [rune(0x1D51B)]
		'xfr;':                             [rune(0x1D535)]
		'xhArr;':                           [rune(0x027FA)]
		'xharr;':                           [rune(0x027F7)]
		'Xi;':                              [rune(0x0039E)]
		'xi;':                              [rune(0x003BE)]
		'xlArr;':                           [rune(0x027F8)]
		'xlarr;':                           [rune(0x027F5)]
		'xmap;':                            [rune(0x027FC)]
		'xnis;':                            [rune(0x022FB)]
		'xodot;':                           [rune(0x02A00)]
		'Xopf;':                            [rune(0x1D54F)]
		'xopf;':                            [rune(0x1D569)]
		'xoplus;':                          [rune(0x02A01)]
		'xotime;':                          [rune(0x02A02)]
		'xrArr;':                           [rune(0x027F9)]
		'xrarr;':                           [rune(0x027F6)]
		'Xscr;':                            [rune(0x1D4B3)]
		'xscr;':                            [rune(0x1D4CD)]
		'xsqcup;':                          [rune(0x02A06)]
		'xuplus;':                          [rune(0x02A04)]
		'xutri;':                           [rune(0x025B3)]
		'xvee;':                            [rune(0x022C1)]
		'xwedge;':                          [rune(0x022C0)]
		'Yacute;':                          [rune(0x000DD)]
		'Yacute':                           [rune(0x000DD)]
		'yacute;':                          [rune(0x000FD)]
		'yacute':                           [rune(0x000FD)]
		'YAcy;':                            [rune(0x0042F)]
		'yacy;':                            [rune(0x0044F)]
		'Ycirc;':                           [rune(0x00176)]
		'ycirc;':                           [rune(0x00177)]
		'Ycy;':                             [rune(0x0042B)]
		'ycy;':                             [rune(0x0044B)]
		'yen;':                             [rune(0x000A5)]
		'yen':                              [rune(0x000A5)]
		'Yfr;':                             [rune(0x1D51C)]
		'yfr;':                             [rune(0x1D536)]
		'YIcy;':                            [rune(0x00407)]
		'yicy;':                            [rune(0x00457)]
		'Yopf;':                            [rune(0x1D550)]
		'yopf;':                            [rune(0x1D56A)]
		'Yscr;':                            [rune(0x1D4B4)]
		'yscr;':                            [rune(0x1D4CE)]
		'YUcy;':                            [rune(0x0042E)]
		'yucy;':                            [rune(0x0044E)]
		'Yuml;':                            [rune(0x00178)]
		'yuml;':                            [rune(0x000FF)]
		'yuml':                             [rune(0x000FF)]
		'Zacute;':                          [rune(0x00179)]
		'zacute;':                          [rune(0x0017A)]
		'Zcaron;':                          [rune(0x0017D)]
		'zcaron;':                          [rune(0x0017E)]
		'Zcy;':                             [rune(0x00417)]
		'zcy;':                             [rune(0x00437)]
		'Zdot;':                            [rune(0x0017B)]
		'zdot;':                            [rune(0x0017C)]
		'zeetrf;':                          [rune(0x02128)]
		'ZeroWidthSpace;':                  [rune(0x0200B)]
		'Zeta;':                            [rune(0x00396)]
		'zeta;':                            [rune(0x003B6)]
		'Zfr;':                             [rune(0x02128)]
		'zfr;':                             [rune(0x1D537)]
		'ZHcy;':                            [rune(0x00416)]
		'zhcy;':                            [rune(0x00436)]
		'zigrarr;':                         [rune(0x021DD)]
		'Zopf;':                            [rune(0x02124)]
		'zopf;':                            [rune(0x1D56B)]
		'Zscr;':                            [rune(0x1D4B5)]
		'zscr;':                            [rune(0x1D4CF)]
		'zwj;':                             [rune(0x0200D)]
		'zwnj;':                            [rune(0x0200C)]
	}
)
