module tokenizer

enum ParseError {
	unexpected_null_character
}