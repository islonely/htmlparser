module htmlparser